magic
tech sky130B
magscale 1 2
timestamp 1666302226
<< nwell >>
rect -858 -40467 858 40467
<< mvpmos >>
rect -600 35370 600 40170
rect -600 30334 600 35134
rect -600 25298 600 30098
rect -600 20262 600 25062
rect -600 15226 600 20026
rect -600 10190 600 14990
rect -600 5154 600 9954
rect -600 118 600 4918
rect -600 -4918 600 -118
rect -600 -9954 600 -5154
rect -600 -14990 600 -10190
rect -600 -20026 600 -15226
rect -600 -25062 600 -20262
rect -600 -30098 600 -25298
rect -600 -35134 600 -30334
rect -600 -40170 600 -35370
<< mvpdiff >>
rect -658 40158 -600 40170
rect -658 35382 -646 40158
rect -612 35382 -600 40158
rect -658 35370 -600 35382
rect 600 40158 658 40170
rect 600 35382 612 40158
rect 646 35382 658 40158
rect 600 35370 658 35382
rect -658 35122 -600 35134
rect -658 30346 -646 35122
rect -612 30346 -600 35122
rect -658 30334 -600 30346
rect 600 35122 658 35134
rect 600 30346 612 35122
rect 646 30346 658 35122
rect 600 30334 658 30346
rect -658 30086 -600 30098
rect -658 25310 -646 30086
rect -612 25310 -600 30086
rect -658 25298 -600 25310
rect 600 30086 658 30098
rect 600 25310 612 30086
rect 646 25310 658 30086
rect 600 25298 658 25310
rect -658 25050 -600 25062
rect -658 20274 -646 25050
rect -612 20274 -600 25050
rect -658 20262 -600 20274
rect 600 25050 658 25062
rect 600 20274 612 25050
rect 646 20274 658 25050
rect 600 20262 658 20274
rect -658 20014 -600 20026
rect -658 15238 -646 20014
rect -612 15238 -600 20014
rect -658 15226 -600 15238
rect 600 20014 658 20026
rect 600 15238 612 20014
rect 646 15238 658 20014
rect 600 15226 658 15238
rect -658 14978 -600 14990
rect -658 10202 -646 14978
rect -612 10202 -600 14978
rect -658 10190 -600 10202
rect 600 14978 658 14990
rect 600 10202 612 14978
rect 646 10202 658 14978
rect 600 10190 658 10202
rect -658 9942 -600 9954
rect -658 5166 -646 9942
rect -612 5166 -600 9942
rect -658 5154 -600 5166
rect 600 9942 658 9954
rect 600 5166 612 9942
rect 646 5166 658 9942
rect 600 5154 658 5166
rect -658 4906 -600 4918
rect -658 130 -646 4906
rect -612 130 -600 4906
rect -658 118 -600 130
rect 600 4906 658 4918
rect 600 130 612 4906
rect 646 130 658 4906
rect 600 118 658 130
rect -658 -130 -600 -118
rect -658 -4906 -646 -130
rect -612 -4906 -600 -130
rect -658 -4918 -600 -4906
rect 600 -130 658 -118
rect 600 -4906 612 -130
rect 646 -4906 658 -130
rect 600 -4918 658 -4906
rect -658 -5166 -600 -5154
rect -658 -9942 -646 -5166
rect -612 -9942 -600 -5166
rect -658 -9954 -600 -9942
rect 600 -5166 658 -5154
rect 600 -9942 612 -5166
rect 646 -9942 658 -5166
rect 600 -9954 658 -9942
rect -658 -10202 -600 -10190
rect -658 -14978 -646 -10202
rect -612 -14978 -600 -10202
rect -658 -14990 -600 -14978
rect 600 -10202 658 -10190
rect 600 -14978 612 -10202
rect 646 -14978 658 -10202
rect 600 -14990 658 -14978
rect -658 -15238 -600 -15226
rect -658 -20014 -646 -15238
rect -612 -20014 -600 -15238
rect -658 -20026 -600 -20014
rect 600 -15238 658 -15226
rect 600 -20014 612 -15238
rect 646 -20014 658 -15238
rect 600 -20026 658 -20014
rect -658 -20274 -600 -20262
rect -658 -25050 -646 -20274
rect -612 -25050 -600 -20274
rect -658 -25062 -600 -25050
rect 600 -20274 658 -20262
rect 600 -25050 612 -20274
rect 646 -25050 658 -20274
rect 600 -25062 658 -25050
rect -658 -25310 -600 -25298
rect -658 -30086 -646 -25310
rect -612 -30086 -600 -25310
rect -658 -30098 -600 -30086
rect 600 -25310 658 -25298
rect 600 -30086 612 -25310
rect 646 -30086 658 -25310
rect 600 -30098 658 -30086
rect -658 -30346 -600 -30334
rect -658 -35122 -646 -30346
rect -612 -35122 -600 -30346
rect -658 -35134 -600 -35122
rect 600 -30346 658 -30334
rect 600 -35122 612 -30346
rect 646 -35122 658 -30346
rect 600 -35134 658 -35122
rect -658 -35382 -600 -35370
rect -658 -40158 -646 -35382
rect -612 -40158 -600 -35382
rect -658 -40170 -600 -40158
rect 600 -35382 658 -35370
rect 600 -40158 612 -35382
rect 646 -40158 658 -35382
rect 600 -40170 658 -40158
<< mvpdiffc >>
rect -646 35382 -612 40158
rect 612 35382 646 40158
rect -646 30346 -612 35122
rect 612 30346 646 35122
rect -646 25310 -612 30086
rect 612 25310 646 30086
rect -646 20274 -612 25050
rect 612 20274 646 25050
rect -646 15238 -612 20014
rect 612 15238 646 20014
rect -646 10202 -612 14978
rect 612 10202 646 14978
rect -646 5166 -612 9942
rect 612 5166 646 9942
rect -646 130 -612 4906
rect 612 130 646 4906
rect -646 -4906 -612 -130
rect 612 -4906 646 -130
rect -646 -9942 -612 -5166
rect 612 -9942 646 -5166
rect -646 -14978 -612 -10202
rect 612 -14978 646 -10202
rect -646 -20014 -612 -15238
rect 612 -20014 646 -15238
rect -646 -25050 -612 -20274
rect 612 -25050 646 -20274
rect -646 -30086 -612 -25310
rect 612 -30086 646 -25310
rect -646 -35122 -612 -30346
rect 612 -35122 646 -30346
rect -646 -40158 -612 -35382
rect 612 -40158 646 -35382
<< mvnsubdiff >>
rect -792 40389 792 40401
rect -792 40355 -684 40389
rect 684 40355 792 40389
rect -792 40343 792 40355
rect -792 40293 -734 40343
rect -792 -40293 -780 40293
rect -746 -40293 -734 40293
rect 734 40293 792 40343
rect -792 -40343 -734 -40293
rect 734 -40293 746 40293
rect 780 -40293 792 40293
rect 734 -40343 792 -40293
rect -792 -40355 792 -40343
rect -792 -40389 -684 -40355
rect 684 -40389 792 -40355
rect -792 -40401 792 -40389
<< mvnsubdiffcont >>
rect -684 40355 684 40389
rect -780 -40293 -746 40293
rect 746 -40293 780 40293
rect -684 -40389 684 -40355
<< poly >>
rect -600 40251 600 40267
rect -600 40217 -584 40251
rect 584 40217 600 40251
rect -600 40170 600 40217
rect -600 35323 600 35370
rect -600 35289 -584 35323
rect 584 35289 600 35323
rect -600 35273 600 35289
rect -600 35215 600 35231
rect -600 35181 -584 35215
rect 584 35181 600 35215
rect -600 35134 600 35181
rect -600 30287 600 30334
rect -600 30253 -584 30287
rect 584 30253 600 30287
rect -600 30237 600 30253
rect -600 30179 600 30195
rect -600 30145 -584 30179
rect 584 30145 600 30179
rect -600 30098 600 30145
rect -600 25251 600 25298
rect -600 25217 -584 25251
rect 584 25217 600 25251
rect -600 25201 600 25217
rect -600 25143 600 25159
rect -600 25109 -584 25143
rect 584 25109 600 25143
rect -600 25062 600 25109
rect -600 20215 600 20262
rect -600 20181 -584 20215
rect 584 20181 600 20215
rect -600 20165 600 20181
rect -600 20107 600 20123
rect -600 20073 -584 20107
rect 584 20073 600 20107
rect -600 20026 600 20073
rect -600 15179 600 15226
rect -600 15145 -584 15179
rect 584 15145 600 15179
rect -600 15129 600 15145
rect -600 15071 600 15087
rect -600 15037 -584 15071
rect 584 15037 600 15071
rect -600 14990 600 15037
rect -600 10143 600 10190
rect -600 10109 -584 10143
rect 584 10109 600 10143
rect -600 10093 600 10109
rect -600 10035 600 10051
rect -600 10001 -584 10035
rect 584 10001 600 10035
rect -600 9954 600 10001
rect -600 5107 600 5154
rect -600 5073 -584 5107
rect 584 5073 600 5107
rect -600 5057 600 5073
rect -600 4999 600 5015
rect -600 4965 -584 4999
rect 584 4965 600 4999
rect -600 4918 600 4965
rect -600 71 600 118
rect -600 37 -584 71
rect 584 37 600 71
rect -600 21 600 37
rect -600 -37 600 -21
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -600 -118 600 -71
rect -600 -4965 600 -4918
rect -600 -4999 -584 -4965
rect 584 -4999 600 -4965
rect -600 -5015 600 -4999
rect -600 -5073 600 -5057
rect -600 -5107 -584 -5073
rect 584 -5107 600 -5073
rect -600 -5154 600 -5107
rect -600 -10001 600 -9954
rect -600 -10035 -584 -10001
rect 584 -10035 600 -10001
rect -600 -10051 600 -10035
rect -600 -10109 600 -10093
rect -600 -10143 -584 -10109
rect 584 -10143 600 -10109
rect -600 -10190 600 -10143
rect -600 -15037 600 -14990
rect -600 -15071 -584 -15037
rect 584 -15071 600 -15037
rect -600 -15087 600 -15071
rect -600 -15145 600 -15129
rect -600 -15179 -584 -15145
rect 584 -15179 600 -15145
rect -600 -15226 600 -15179
rect -600 -20073 600 -20026
rect -600 -20107 -584 -20073
rect 584 -20107 600 -20073
rect -600 -20123 600 -20107
rect -600 -20181 600 -20165
rect -600 -20215 -584 -20181
rect 584 -20215 600 -20181
rect -600 -20262 600 -20215
rect -600 -25109 600 -25062
rect -600 -25143 -584 -25109
rect 584 -25143 600 -25109
rect -600 -25159 600 -25143
rect -600 -25217 600 -25201
rect -600 -25251 -584 -25217
rect 584 -25251 600 -25217
rect -600 -25298 600 -25251
rect -600 -30145 600 -30098
rect -600 -30179 -584 -30145
rect 584 -30179 600 -30145
rect -600 -30195 600 -30179
rect -600 -30253 600 -30237
rect -600 -30287 -584 -30253
rect 584 -30287 600 -30253
rect -600 -30334 600 -30287
rect -600 -35181 600 -35134
rect -600 -35215 -584 -35181
rect 584 -35215 600 -35181
rect -600 -35231 600 -35215
rect -600 -35289 600 -35273
rect -600 -35323 -584 -35289
rect 584 -35323 600 -35289
rect -600 -35370 600 -35323
rect -600 -40217 600 -40170
rect -600 -40251 -584 -40217
rect 584 -40251 600 -40217
rect -600 -40267 600 -40251
<< polycont >>
rect -584 40217 584 40251
rect -584 35289 584 35323
rect -584 35181 584 35215
rect -584 30253 584 30287
rect -584 30145 584 30179
rect -584 25217 584 25251
rect -584 25109 584 25143
rect -584 20181 584 20215
rect -584 20073 584 20107
rect -584 15145 584 15179
rect -584 15037 584 15071
rect -584 10109 584 10143
rect -584 10001 584 10035
rect -584 5073 584 5107
rect -584 4965 584 4999
rect -584 37 584 71
rect -584 -71 584 -37
rect -584 -4999 584 -4965
rect -584 -5107 584 -5073
rect -584 -10035 584 -10001
rect -584 -10143 584 -10109
rect -584 -15071 584 -15037
rect -584 -15179 584 -15145
rect -584 -20107 584 -20073
rect -584 -20215 584 -20181
rect -584 -25143 584 -25109
rect -584 -25251 584 -25217
rect -584 -30179 584 -30145
rect -584 -30287 584 -30253
rect -584 -35215 584 -35181
rect -584 -35323 584 -35289
rect -584 -40251 584 -40217
<< locali >>
rect -780 40355 -684 40389
rect 684 40355 780 40389
rect -780 40293 -746 40355
rect 746 40293 780 40355
rect -600 40217 -584 40251
rect 584 40217 600 40251
rect -646 40158 -612 40174
rect -646 35366 -612 35382
rect 612 40158 646 40174
rect 612 35366 646 35382
rect -600 35289 -584 35323
rect 584 35289 600 35323
rect -600 35181 -584 35215
rect 584 35181 600 35215
rect -646 35122 -612 35138
rect -646 30330 -612 30346
rect 612 35122 646 35138
rect 612 30330 646 30346
rect -600 30253 -584 30287
rect 584 30253 600 30287
rect -600 30145 -584 30179
rect 584 30145 600 30179
rect -646 30086 -612 30102
rect -646 25294 -612 25310
rect 612 30086 646 30102
rect 612 25294 646 25310
rect -600 25217 -584 25251
rect 584 25217 600 25251
rect -600 25109 -584 25143
rect 584 25109 600 25143
rect -646 25050 -612 25066
rect -646 20258 -612 20274
rect 612 25050 646 25066
rect 612 20258 646 20274
rect -600 20181 -584 20215
rect 584 20181 600 20215
rect -600 20073 -584 20107
rect 584 20073 600 20107
rect -646 20014 -612 20030
rect -646 15222 -612 15238
rect 612 20014 646 20030
rect 612 15222 646 15238
rect -600 15145 -584 15179
rect 584 15145 600 15179
rect -600 15037 -584 15071
rect 584 15037 600 15071
rect -646 14978 -612 14994
rect -646 10186 -612 10202
rect 612 14978 646 14994
rect 612 10186 646 10202
rect -600 10109 -584 10143
rect 584 10109 600 10143
rect -600 10001 -584 10035
rect 584 10001 600 10035
rect -646 9942 -612 9958
rect -646 5150 -612 5166
rect 612 9942 646 9958
rect 612 5150 646 5166
rect -600 5073 -584 5107
rect 584 5073 600 5107
rect -600 4965 -584 4999
rect 584 4965 600 4999
rect -646 4906 -612 4922
rect -646 114 -612 130
rect 612 4906 646 4922
rect 612 114 646 130
rect -600 37 -584 71
rect 584 37 600 71
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -646 -130 -612 -114
rect -646 -4922 -612 -4906
rect 612 -130 646 -114
rect 612 -4922 646 -4906
rect -600 -4999 -584 -4965
rect 584 -4999 600 -4965
rect -600 -5107 -584 -5073
rect 584 -5107 600 -5073
rect -646 -5166 -612 -5150
rect -646 -9958 -612 -9942
rect 612 -5166 646 -5150
rect 612 -9958 646 -9942
rect -600 -10035 -584 -10001
rect 584 -10035 600 -10001
rect -600 -10143 -584 -10109
rect 584 -10143 600 -10109
rect -646 -10202 -612 -10186
rect -646 -14994 -612 -14978
rect 612 -10202 646 -10186
rect 612 -14994 646 -14978
rect -600 -15071 -584 -15037
rect 584 -15071 600 -15037
rect -600 -15179 -584 -15145
rect 584 -15179 600 -15145
rect -646 -15238 -612 -15222
rect -646 -20030 -612 -20014
rect 612 -15238 646 -15222
rect 612 -20030 646 -20014
rect -600 -20107 -584 -20073
rect 584 -20107 600 -20073
rect -600 -20215 -584 -20181
rect 584 -20215 600 -20181
rect -646 -20274 -612 -20258
rect -646 -25066 -612 -25050
rect 612 -20274 646 -20258
rect 612 -25066 646 -25050
rect -600 -25143 -584 -25109
rect 584 -25143 600 -25109
rect -600 -25251 -584 -25217
rect 584 -25251 600 -25217
rect -646 -25310 -612 -25294
rect -646 -30102 -612 -30086
rect 612 -25310 646 -25294
rect 612 -30102 646 -30086
rect -600 -30179 -584 -30145
rect 584 -30179 600 -30145
rect -600 -30287 -584 -30253
rect 584 -30287 600 -30253
rect -646 -30346 -612 -30330
rect -646 -35138 -612 -35122
rect 612 -30346 646 -30330
rect 612 -35138 646 -35122
rect -600 -35215 -584 -35181
rect 584 -35215 600 -35181
rect -600 -35323 -584 -35289
rect 584 -35323 600 -35289
rect -646 -35382 -612 -35366
rect -646 -40174 -612 -40158
rect 612 -35382 646 -35366
rect 612 -40174 646 -40158
rect -600 -40251 -584 -40217
rect 584 -40251 600 -40217
rect -780 -40355 -746 -40293
rect 746 -40355 780 -40293
rect -780 -40389 -684 -40355
rect 684 -40389 780 -40355
<< viali >>
rect -584 40217 584 40251
rect -646 35382 -612 40158
rect 612 35382 646 40158
rect -584 35289 584 35323
rect -584 35181 584 35215
rect -646 30346 -612 35122
rect 612 30346 646 35122
rect -584 30253 584 30287
rect -584 30145 584 30179
rect -646 25310 -612 30086
rect 612 25310 646 30086
rect -584 25217 584 25251
rect -584 25109 584 25143
rect -646 20274 -612 25050
rect 612 20274 646 25050
rect -584 20181 584 20215
rect -584 20073 584 20107
rect -646 15238 -612 20014
rect 612 15238 646 20014
rect -584 15145 584 15179
rect -584 15037 584 15071
rect -646 10202 -612 14978
rect 612 10202 646 14978
rect -584 10109 584 10143
rect -584 10001 584 10035
rect -646 5166 -612 9942
rect 612 5166 646 9942
rect -584 5073 584 5107
rect -584 4965 584 4999
rect -646 130 -612 4906
rect 612 130 646 4906
rect -584 37 584 71
rect -584 -71 584 -37
rect -646 -4906 -612 -130
rect 612 -4906 646 -130
rect -584 -4999 584 -4965
rect -584 -5107 584 -5073
rect -646 -9942 -612 -5166
rect 612 -9942 646 -5166
rect -584 -10035 584 -10001
rect -584 -10143 584 -10109
rect -646 -14978 -612 -10202
rect 612 -14978 646 -10202
rect -584 -15071 584 -15037
rect -584 -15179 584 -15145
rect -646 -20014 -612 -15238
rect 612 -20014 646 -15238
rect -584 -20107 584 -20073
rect -584 -20215 584 -20181
rect -646 -25050 -612 -20274
rect 612 -25050 646 -20274
rect -584 -25143 584 -25109
rect -584 -25251 584 -25217
rect -646 -30086 -612 -25310
rect 612 -30086 646 -25310
rect -584 -30179 584 -30145
rect -584 -30287 584 -30253
rect -646 -35122 -612 -30346
rect 612 -35122 646 -30346
rect -584 -35215 584 -35181
rect -584 -35323 584 -35289
rect -646 -40158 -612 -35382
rect 612 -40158 646 -35382
rect -584 -40251 584 -40217
<< metal1 >>
rect -596 40251 596 40257
rect -596 40217 -584 40251
rect 584 40217 596 40251
rect -596 40211 596 40217
rect -652 40158 -606 40170
rect -652 35382 -646 40158
rect -612 35382 -606 40158
rect -652 35370 -606 35382
rect 606 40158 652 40170
rect 606 35382 612 40158
rect 646 35382 652 40158
rect 606 35370 652 35382
rect -596 35323 596 35329
rect -596 35289 -584 35323
rect 584 35289 596 35323
rect -596 35283 596 35289
rect -596 35215 596 35221
rect -596 35181 -584 35215
rect 584 35181 596 35215
rect -596 35175 596 35181
rect -652 35122 -606 35134
rect -652 30346 -646 35122
rect -612 30346 -606 35122
rect -652 30334 -606 30346
rect 606 35122 652 35134
rect 606 30346 612 35122
rect 646 30346 652 35122
rect 606 30334 652 30346
rect -596 30287 596 30293
rect -596 30253 -584 30287
rect 584 30253 596 30287
rect -596 30247 596 30253
rect -596 30179 596 30185
rect -596 30145 -584 30179
rect 584 30145 596 30179
rect -596 30139 596 30145
rect -652 30086 -606 30098
rect -652 25310 -646 30086
rect -612 25310 -606 30086
rect -652 25298 -606 25310
rect 606 30086 652 30098
rect 606 25310 612 30086
rect 646 25310 652 30086
rect 606 25298 652 25310
rect -596 25251 596 25257
rect -596 25217 -584 25251
rect 584 25217 596 25251
rect -596 25211 596 25217
rect -596 25143 596 25149
rect -596 25109 -584 25143
rect 584 25109 596 25143
rect -596 25103 596 25109
rect -652 25050 -606 25062
rect -652 20274 -646 25050
rect -612 20274 -606 25050
rect -652 20262 -606 20274
rect 606 25050 652 25062
rect 606 20274 612 25050
rect 646 20274 652 25050
rect 606 20262 652 20274
rect -596 20215 596 20221
rect -596 20181 -584 20215
rect 584 20181 596 20215
rect -596 20175 596 20181
rect -596 20107 596 20113
rect -596 20073 -584 20107
rect 584 20073 596 20107
rect -596 20067 596 20073
rect -652 20014 -606 20026
rect -652 15238 -646 20014
rect -612 15238 -606 20014
rect -652 15226 -606 15238
rect 606 20014 652 20026
rect 606 15238 612 20014
rect 646 15238 652 20014
rect 606 15226 652 15238
rect -596 15179 596 15185
rect -596 15145 -584 15179
rect 584 15145 596 15179
rect -596 15139 596 15145
rect -596 15071 596 15077
rect -596 15037 -584 15071
rect 584 15037 596 15071
rect -596 15031 596 15037
rect -652 14978 -606 14990
rect -652 10202 -646 14978
rect -612 10202 -606 14978
rect -652 10190 -606 10202
rect 606 14978 652 14990
rect 606 10202 612 14978
rect 646 10202 652 14978
rect 606 10190 652 10202
rect -596 10143 596 10149
rect -596 10109 -584 10143
rect 584 10109 596 10143
rect -596 10103 596 10109
rect -596 10035 596 10041
rect -596 10001 -584 10035
rect 584 10001 596 10035
rect -596 9995 596 10001
rect -652 9942 -606 9954
rect -652 5166 -646 9942
rect -612 5166 -606 9942
rect -652 5154 -606 5166
rect 606 9942 652 9954
rect 606 5166 612 9942
rect 646 5166 652 9942
rect 606 5154 652 5166
rect -596 5107 596 5113
rect -596 5073 -584 5107
rect 584 5073 596 5107
rect -596 5067 596 5073
rect -596 4999 596 5005
rect -596 4965 -584 4999
rect 584 4965 596 4999
rect -596 4959 596 4965
rect -652 4906 -606 4918
rect -652 130 -646 4906
rect -612 130 -606 4906
rect -652 118 -606 130
rect 606 4906 652 4918
rect 606 130 612 4906
rect 646 130 652 4906
rect 606 118 652 130
rect -596 71 596 77
rect -596 37 -584 71
rect 584 37 596 71
rect -596 31 596 37
rect -596 -37 596 -31
rect -596 -71 -584 -37
rect 584 -71 596 -37
rect -596 -77 596 -71
rect -652 -130 -606 -118
rect -652 -4906 -646 -130
rect -612 -4906 -606 -130
rect -652 -4918 -606 -4906
rect 606 -130 652 -118
rect 606 -4906 612 -130
rect 646 -4906 652 -130
rect 606 -4918 652 -4906
rect -596 -4965 596 -4959
rect -596 -4999 -584 -4965
rect 584 -4999 596 -4965
rect -596 -5005 596 -4999
rect -596 -5073 596 -5067
rect -596 -5107 -584 -5073
rect 584 -5107 596 -5073
rect -596 -5113 596 -5107
rect -652 -5166 -606 -5154
rect -652 -9942 -646 -5166
rect -612 -9942 -606 -5166
rect -652 -9954 -606 -9942
rect 606 -5166 652 -5154
rect 606 -9942 612 -5166
rect 646 -9942 652 -5166
rect 606 -9954 652 -9942
rect -596 -10001 596 -9995
rect -596 -10035 -584 -10001
rect 584 -10035 596 -10001
rect -596 -10041 596 -10035
rect -596 -10109 596 -10103
rect -596 -10143 -584 -10109
rect 584 -10143 596 -10109
rect -596 -10149 596 -10143
rect -652 -10202 -606 -10190
rect -652 -14978 -646 -10202
rect -612 -14978 -606 -10202
rect -652 -14990 -606 -14978
rect 606 -10202 652 -10190
rect 606 -14978 612 -10202
rect 646 -14978 652 -10202
rect 606 -14990 652 -14978
rect -596 -15037 596 -15031
rect -596 -15071 -584 -15037
rect 584 -15071 596 -15037
rect -596 -15077 596 -15071
rect -596 -15145 596 -15139
rect -596 -15179 -584 -15145
rect 584 -15179 596 -15145
rect -596 -15185 596 -15179
rect -652 -15238 -606 -15226
rect -652 -20014 -646 -15238
rect -612 -20014 -606 -15238
rect -652 -20026 -606 -20014
rect 606 -15238 652 -15226
rect 606 -20014 612 -15238
rect 646 -20014 652 -15238
rect 606 -20026 652 -20014
rect -596 -20073 596 -20067
rect -596 -20107 -584 -20073
rect 584 -20107 596 -20073
rect -596 -20113 596 -20107
rect -596 -20181 596 -20175
rect -596 -20215 -584 -20181
rect 584 -20215 596 -20181
rect -596 -20221 596 -20215
rect -652 -20274 -606 -20262
rect -652 -25050 -646 -20274
rect -612 -25050 -606 -20274
rect -652 -25062 -606 -25050
rect 606 -20274 652 -20262
rect 606 -25050 612 -20274
rect 646 -25050 652 -20274
rect 606 -25062 652 -25050
rect -596 -25109 596 -25103
rect -596 -25143 -584 -25109
rect 584 -25143 596 -25109
rect -596 -25149 596 -25143
rect -596 -25217 596 -25211
rect -596 -25251 -584 -25217
rect 584 -25251 596 -25217
rect -596 -25257 596 -25251
rect -652 -25310 -606 -25298
rect -652 -30086 -646 -25310
rect -612 -30086 -606 -25310
rect -652 -30098 -606 -30086
rect 606 -25310 652 -25298
rect 606 -30086 612 -25310
rect 646 -30086 652 -25310
rect 606 -30098 652 -30086
rect -596 -30145 596 -30139
rect -596 -30179 -584 -30145
rect 584 -30179 596 -30145
rect -596 -30185 596 -30179
rect -596 -30253 596 -30247
rect -596 -30287 -584 -30253
rect 584 -30287 596 -30253
rect -596 -30293 596 -30287
rect -652 -30346 -606 -30334
rect -652 -35122 -646 -30346
rect -612 -35122 -606 -30346
rect -652 -35134 -606 -35122
rect 606 -30346 652 -30334
rect 606 -35122 612 -30346
rect 646 -35122 652 -30346
rect 606 -35134 652 -35122
rect -596 -35181 596 -35175
rect -596 -35215 -584 -35181
rect 584 -35215 596 -35181
rect -596 -35221 596 -35215
rect -596 -35289 596 -35283
rect -596 -35323 -584 -35289
rect 584 -35323 596 -35289
rect -596 -35329 596 -35323
rect -652 -35382 -606 -35370
rect -652 -40158 -646 -35382
rect -612 -40158 -606 -35382
rect -652 -40170 -606 -40158
rect 606 -35382 652 -35370
rect 606 -40158 612 -35382
rect 646 -40158 652 -35382
rect 606 -40170 652 -40158
rect -596 -40217 596 -40211
rect -596 -40251 -584 -40217
rect 584 -40251 596 -40217
rect -596 -40257 596 -40251
<< properties >>
string FIXED_BBOX -763 -40372 763 40372
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 24.0 l 6.0 m 16 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
