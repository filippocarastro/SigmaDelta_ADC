magic
tech sky130B
magscale 1 2
timestamp 1667934541
<< error_p >>
rect -3240 3298 3240 3302
rect -3240 -3230 -3210 3298
rect -3174 3232 3174 3236
rect -3174 -3164 -3144 3232
rect 3144 -3164 3174 3232
rect 3210 -3230 3240 3298
<< nwell >>
rect -3210 -3264 3210 3298
<< mvpmos >>
rect -3116 -3164 -1916 3236
rect -1858 -3164 -658 3236
rect -600 -3164 600 3236
rect 658 -3164 1858 3236
rect 1916 -3164 3116 3236
<< mvpdiff >>
rect -3174 2586 -3116 3236
rect -3174 -2514 -3162 2586
rect -3128 -2514 -3116 2586
rect -3174 -3164 -3116 -2514
rect -1916 2586 -1858 3236
rect -1916 -2514 -1904 2586
rect -1870 -2514 -1858 2586
rect -1916 -3164 -1858 -2514
rect -658 2586 -600 3236
rect -658 -2514 -646 2586
rect -612 -2514 -600 2586
rect -658 -3164 -600 -2514
rect 600 2586 658 3236
rect 600 -2514 612 2586
rect 646 -2514 658 2586
rect 600 -3164 658 -2514
rect 1858 2586 1916 3236
rect 1858 -2514 1870 2586
rect 1904 -2514 1916 2586
rect 1858 -3164 1916 -2514
rect 3116 2586 3174 3236
rect 3116 -2514 3128 2586
rect 3162 -2514 3174 2586
rect 3116 -3164 3174 -2514
<< mvpdiffc >>
rect -3162 -2514 -3128 2586
rect -1904 -2514 -1870 2586
rect -646 -2514 -612 2586
rect 612 -2514 646 2586
rect 1870 -2514 1904 2586
rect 3128 -2514 3162 2586
<< poly >>
rect -3116 3236 -1916 3262
rect -1858 3236 -658 3262
rect -600 3236 600 3262
rect 658 3236 1858 3262
rect 1916 3236 3116 3262
rect -3116 -3211 -1916 -3164
rect -3116 -3228 -3042 -3211
rect -3058 -3245 -3042 -3228
rect -1990 -3228 -1916 -3211
rect -1858 -3211 -658 -3164
rect -1858 -3228 -1784 -3211
rect -1990 -3245 -1974 -3228
rect -3058 -3261 -1974 -3245
rect -1800 -3245 -1784 -3228
rect -732 -3228 -658 -3211
rect -600 -3211 600 -3164
rect -600 -3228 -526 -3211
rect -732 -3245 -716 -3228
rect -1800 -3261 -716 -3245
rect -542 -3245 -526 -3228
rect 526 -3228 600 -3211
rect 658 -3211 1858 -3164
rect 658 -3228 732 -3211
rect 526 -3245 542 -3228
rect -542 -3261 542 -3245
rect 716 -3245 732 -3228
rect 1784 -3228 1858 -3211
rect 1916 -3211 3116 -3164
rect 1916 -3228 1990 -3211
rect 1784 -3245 1800 -3228
rect 716 -3261 1800 -3245
rect 1974 -3245 1990 -3228
rect 3042 -3228 3116 -3211
rect 3042 -3245 3058 -3228
rect 1974 -3261 3058 -3245
<< polycont >>
rect -3042 -3245 -1990 -3211
rect -1784 -3245 -732 -3211
rect -526 -3245 526 -3211
rect 732 -3245 1784 -3211
rect 1990 -3245 3042 -3211
<< locali >>
rect -3162 2586 -3128 2602
rect -3162 -2530 -3128 -2514
rect -1904 2586 -1870 2602
rect -1904 -2530 -1870 -2514
rect -646 2586 -612 2602
rect -646 -2530 -612 -2514
rect 612 2586 646 2602
rect 612 -2530 646 -2514
rect 1870 2586 1904 2602
rect 1870 -2530 1904 -2514
rect 3128 2586 3162 2602
rect 3128 -2530 3162 -2514
rect -3058 -3245 -3042 -3211
rect -1990 -3245 -1974 -3211
rect -1800 -3245 -1784 -3211
rect -732 -3245 -716 -3211
rect -542 -3245 -526 -3211
rect 526 -3245 542 -3211
rect 716 -3245 732 -3211
rect 1784 -3245 1800 -3211
rect 1974 -3245 1990 -3211
rect 3042 -3245 3058 -3211
<< viali >>
rect -3162 -2514 -3128 2586
rect -1904 -2514 -1870 2586
rect -646 -2514 -612 2586
rect 612 -2514 646 2586
rect 1870 -2514 1904 2586
rect 3128 -2514 3162 2586
rect -3042 -3245 -1990 -3211
rect -1784 -3245 -732 -3211
rect -526 -3245 526 -3211
rect 732 -3245 1784 -3211
rect 1990 -3245 3042 -3211
<< metal1 >>
rect -3168 2586 -3122 2598
rect -3168 -2514 -3162 2586
rect -3128 -2514 -3122 2586
rect -3168 -2526 -3122 -2514
rect -1910 2586 -1864 2598
rect -1910 -2514 -1904 2586
rect -1870 -2514 -1864 2586
rect -1910 -2526 -1864 -2514
rect -652 2586 -606 2598
rect -652 -2514 -646 2586
rect -612 -2514 -606 2586
rect -652 -2526 -606 -2514
rect 606 2586 652 2598
rect 606 -2514 612 2586
rect 646 -2514 652 2586
rect 606 -2526 652 -2514
rect 1864 2586 1910 2598
rect 1864 -2514 1870 2586
rect 1904 -2514 1910 2586
rect 1864 -2526 1910 -2514
rect 3122 2586 3168 2598
rect 3122 -2514 3128 2586
rect 3162 -2514 3168 2586
rect 3122 -2526 3168 -2514
rect -3054 -3211 -1978 -3205
rect -3054 -3245 -3042 -3211
rect -1990 -3245 -1978 -3211
rect -3054 -3251 -1978 -3245
rect -1796 -3211 -720 -3205
rect -1796 -3245 -1784 -3211
rect -732 -3245 -720 -3211
rect -1796 -3251 -720 -3245
rect -538 -3211 538 -3205
rect -538 -3245 -526 -3211
rect 526 -3245 538 -3211
rect -538 -3251 538 -3245
rect 720 -3211 1796 -3205
rect 720 -3245 732 -3211
rect 1784 -3245 1796 -3211
rect 720 -3251 1796 -3245
rect 1978 -3211 3054 -3205
rect 1978 -3245 1990 -3211
rect 3042 -3245 3054 -3211
rect 1978 -3251 3054 -3245
<< properties >>
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 6.0 m 1 nf 5 diffcov 80 polycov 90 guard 0 glc 0 grc 0 gtc 0 gbc 0 tbcov 80 rlcov 80 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 80 viadrn 80 viagate 90 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
