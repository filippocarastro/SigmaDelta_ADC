magic
tech sky130B
magscale 1 2
timestamp 1667069721
<< nwell >>
rect -10293 -2697 10293 2697
<< mvpmos >>
rect -10035 -2400 -8835 2400
rect -8777 -2400 -7577 2400
rect -7519 -2400 -6319 2400
rect -6261 -2400 -5061 2400
rect -5003 -2400 -3803 2400
rect -3745 -2400 -2545 2400
rect -2487 -2400 -1287 2400
rect -1229 -2400 -29 2400
rect 29 -2400 1229 2400
rect 1287 -2400 2487 2400
rect 2545 -2400 3745 2400
rect 3803 -2400 5003 2400
rect 5061 -2400 6261 2400
rect 6319 -2400 7519 2400
rect 7577 -2400 8777 2400
rect 8835 -2400 10035 2400
<< mvpdiff >>
rect -10093 2388 -10035 2400
rect -10093 -2388 -10081 2388
rect -10047 -2388 -10035 2388
rect -10093 -2400 -10035 -2388
rect -8835 2388 -8777 2400
rect -8835 -2388 -8823 2388
rect -8789 -2388 -8777 2388
rect -8835 -2400 -8777 -2388
rect -7577 2388 -7519 2400
rect -7577 -2388 -7565 2388
rect -7531 -2388 -7519 2388
rect -7577 -2400 -7519 -2388
rect -6319 2388 -6261 2400
rect -6319 -2388 -6307 2388
rect -6273 -2388 -6261 2388
rect -6319 -2400 -6261 -2388
rect -5061 2388 -5003 2400
rect -5061 -2388 -5049 2388
rect -5015 -2388 -5003 2388
rect -5061 -2400 -5003 -2388
rect -3803 2388 -3745 2400
rect -3803 -2388 -3791 2388
rect -3757 -2388 -3745 2388
rect -3803 -2400 -3745 -2388
rect -2545 2388 -2487 2400
rect -2545 -2388 -2533 2388
rect -2499 -2388 -2487 2388
rect -2545 -2400 -2487 -2388
rect -1287 2388 -1229 2400
rect -1287 -2388 -1275 2388
rect -1241 -2388 -1229 2388
rect -1287 -2400 -1229 -2388
rect -29 2388 29 2400
rect -29 -2388 -17 2388
rect 17 -2388 29 2388
rect -29 -2400 29 -2388
rect 1229 2388 1287 2400
rect 1229 -2388 1241 2388
rect 1275 -2388 1287 2388
rect 1229 -2400 1287 -2388
rect 2487 2388 2545 2400
rect 2487 -2388 2499 2388
rect 2533 -2388 2545 2388
rect 2487 -2400 2545 -2388
rect 3745 2388 3803 2400
rect 3745 -2388 3757 2388
rect 3791 -2388 3803 2388
rect 3745 -2400 3803 -2388
rect 5003 2388 5061 2400
rect 5003 -2388 5015 2388
rect 5049 -2388 5061 2388
rect 5003 -2400 5061 -2388
rect 6261 2388 6319 2400
rect 6261 -2388 6273 2388
rect 6307 -2388 6319 2388
rect 6261 -2400 6319 -2388
rect 7519 2388 7577 2400
rect 7519 -2388 7531 2388
rect 7565 -2388 7577 2388
rect 7519 -2400 7577 -2388
rect 8777 2388 8835 2400
rect 8777 -2388 8789 2388
rect 8823 -2388 8835 2388
rect 8777 -2400 8835 -2388
rect 10035 2388 10093 2400
rect 10035 -2388 10047 2388
rect 10081 -2388 10093 2388
rect 10035 -2400 10093 -2388
<< mvpdiffc >>
rect -10081 -2388 -10047 2388
rect -8823 -2388 -8789 2388
rect -7565 -2388 -7531 2388
rect -6307 -2388 -6273 2388
rect -5049 -2388 -5015 2388
rect -3791 -2388 -3757 2388
rect -2533 -2388 -2499 2388
rect -1275 -2388 -1241 2388
rect -17 -2388 17 2388
rect 1241 -2388 1275 2388
rect 2499 -2388 2533 2388
rect 3757 -2388 3791 2388
rect 5015 -2388 5049 2388
rect 6273 -2388 6307 2388
rect 7531 -2388 7565 2388
rect 8789 -2388 8823 2388
rect 10047 -2388 10081 2388
<< mvnsubdiff >>
rect -10227 2619 10227 2631
rect -10227 2585 -10119 2619
rect 10119 2585 10227 2619
rect -10227 2573 10227 2585
rect -10227 2523 -10169 2573
rect -10227 -2523 -10215 2523
rect -10181 -2523 -10169 2523
rect 10169 2523 10227 2573
rect -10227 -2573 -10169 -2523
rect 10169 -2523 10181 2523
rect 10215 -2523 10227 2523
rect 10169 -2573 10227 -2523
rect -10227 -2585 10227 -2573
rect -10227 -2619 -10119 -2585
rect 10119 -2619 10227 -2585
rect -10227 -2631 10227 -2619
<< mvnsubdiffcont >>
rect -10119 2585 10119 2619
rect -10215 -2523 -10181 2523
rect 10181 -2523 10215 2523
rect -10119 -2619 10119 -2585
<< poly >>
rect -10035 2481 -8835 2497
rect -10035 2447 -10019 2481
rect -8851 2447 -8835 2481
rect -10035 2400 -8835 2447
rect -8777 2481 -7577 2497
rect -8777 2447 -8761 2481
rect -7593 2447 -7577 2481
rect -8777 2400 -7577 2447
rect -7519 2481 -6319 2497
rect -7519 2447 -7503 2481
rect -6335 2447 -6319 2481
rect -7519 2400 -6319 2447
rect -6261 2481 -5061 2497
rect -6261 2447 -6245 2481
rect -5077 2447 -5061 2481
rect -6261 2400 -5061 2447
rect -5003 2481 -3803 2497
rect -5003 2447 -4987 2481
rect -3819 2447 -3803 2481
rect -5003 2400 -3803 2447
rect -3745 2481 -2545 2497
rect -3745 2447 -3729 2481
rect -2561 2447 -2545 2481
rect -3745 2400 -2545 2447
rect -2487 2481 -1287 2497
rect -2487 2447 -2471 2481
rect -1303 2447 -1287 2481
rect -2487 2400 -1287 2447
rect -1229 2481 -29 2497
rect -1229 2447 -1213 2481
rect -45 2447 -29 2481
rect -1229 2400 -29 2447
rect 29 2481 1229 2497
rect 29 2447 45 2481
rect 1213 2447 1229 2481
rect 29 2400 1229 2447
rect 1287 2481 2487 2497
rect 1287 2447 1303 2481
rect 2471 2447 2487 2481
rect 1287 2400 2487 2447
rect 2545 2481 3745 2497
rect 2545 2447 2561 2481
rect 3729 2447 3745 2481
rect 2545 2400 3745 2447
rect 3803 2481 5003 2497
rect 3803 2447 3819 2481
rect 4987 2447 5003 2481
rect 3803 2400 5003 2447
rect 5061 2481 6261 2497
rect 5061 2447 5077 2481
rect 6245 2447 6261 2481
rect 5061 2400 6261 2447
rect 6319 2481 7519 2497
rect 6319 2447 6335 2481
rect 7503 2447 7519 2481
rect 6319 2400 7519 2447
rect 7577 2481 8777 2497
rect 7577 2447 7593 2481
rect 8761 2447 8777 2481
rect 7577 2400 8777 2447
rect 8835 2481 10035 2497
rect 8835 2447 8851 2481
rect 10019 2447 10035 2481
rect 8835 2400 10035 2447
rect -10035 -2447 -8835 -2400
rect -10035 -2481 -10019 -2447
rect -8851 -2481 -8835 -2447
rect -10035 -2497 -8835 -2481
rect -8777 -2447 -7577 -2400
rect -8777 -2481 -8761 -2447
rect -7593 -2481 -7577 -2447
rect -8777 -2497 -7577 -2481
rect -7519 -2447 -6319 -2400
rect -7519 -2481 -7503 -2447
rect -6335 -2481 -6319 -2447
rect -7519 -2497 -6319 -2481
rect -6261 -2447 -5061 -2400
rect -6261 -2481 -6245 -2447
rect -5077 -2481 -5061 -2447
rect -6261 -2497 -5061 -2481
rect -5003 -2447 -3803 -2400
rect -5003 -2481 -4987 -2447
rect -3819 -2481 -3803 -2447
rect -5003 -2497 -3803 -2481
rect -3745 -2447 -2545 -2400
rect -3745 -2481 -3729 -2447
rect -2561 -2481 -2545 -2447
rect -3745 -2497 -2545 -2481
rect -2487 -2447 -1287 -2400
rect -2487 -2481 -2471 -2447
rect -1303 -2481 -1287 -2447
rect -2487 -2497 -1287 -2481
rect -1229 -2447 -29 -2400
rect -1229 -2481 -1213 -2447
rect -45 -2481 -29 -2447
rect -1229 -2497 -29 -2481
rect 29 -2447 1229 -2400
rect 29 -2481 45 -2447
rect 1213 -2481 1229 -2447
rect 29 -2497 1229 -2481
rect 1287 -2447 2487 -2400
rect 1287 -2481 1303 -2447
rect 2471 -2481 2487 -2447
rect 1287 -2497 2487 -2481
rect 2545 -2447 3745 -2400
rect 2545 -2481 2561 -2447
rect 3729 -2481 3745 -2447
rect 2545 -2497 3745 -2481
rect 3803 -2447 5003 -2400
rect 3803 -2481 3819 -2447
rect 4987 -2481 5003 -2447
rect 3803 -2497 5003 -2481
rect 5061 -2447 6261 -2400
rect 5061 -2481 5077 -2447
rect 6245 -2481 6261 -2447
rect 5061 -2497 6261 -2481
rect 6319 -2447 7519 -2400
rect 6319 -2481 6335 -2447
rect 7503 -2481 7519 -2447
rect 6319 -2497 7519 -2481
rect 7577 -2447 8777 -2400
rect 7577 -2481 7593 -2447
rect 8761 -2481 8777 -2447
rect 7577 -2497 8777 -2481
rect 8835 -2447 10035 -2400
rect 8835 -2481 8851 -2447
rect 10019 -2481 10035 -2447
rect 8835 -2497 10035 -2481
<< polycont >>
rect -10019 2447 -8851 2481
rect -8761 2447 -7593 2481
rect -7503 2447 -6335 2481
rect -6245 2447 -5077 2481
rect -4987 2447 -3819 2481
rect -3729 2447 -2561 2481
rect -2471 2447 -1303 2481
rect -1213 2447 -45 2481
rect 45 2447 1213 2481
rect 1303 2447 2471 2481
rect 2561 2447 3729 2481
rect 3819 2447 4987 2481
rect 5077 2447 6245 2481
rect 6335 2447 7503 2481
rect 7593 2447 8761 2481
rect 8851 2447 10019 2481
rect -10019 -2481 -8851 -2447
rect -8761 -2481 -7593 -2447
rect -7503 -2481 -6335 -2447
rect -6245 -2481 -5077 -2447
rect -4987 -2481 -3819 -2447
rect -3729 -2481 -2561 -2447
rect -2471 -2481 -1303 -2447
rect -1213 -2481 -45 -2447
rect 45 -2481 1213 -2447
rect 1303 -2481 2471 -2447
rect 2561 -2481 3729 -2447
rect 3819 -2481 4987 -2447
rect 5077 -2481 6245 -2447
rect 6335 -2481 7503 -2447
rect 7593 -2481 8761 -2447
rect 8851 -2481 10019 -2447
<< locali >>
rect -10215 2585 -10119 2619
rect 10119 2585 10215 2619
rect -10215 2523 -10181 2585
rect 10181 2523 10215 2585
rect -10035 2447 -10019 2481
rect -8851 2447 -8835 2481
rect -8777 2447 -8761 2481
rect -7593 2447 -7577 2481
rect -7519 2447 -7503 2481
rect -6335 2447 -6319 2481
rect -6261 2447 -6245 2481
rect -5077 2447 -5061 2481
rect -5003 2447 -4987 2481
rect -3819 2447 -3803 2481
rect -3745 2447 -3729 2481
rect -2561 2447 -2545 2481
rect -2487 2447 -2471 2481
rect -1303 2447 -1287 2481
rect -1229 2447 -1213 2481
rect -45 2447 -29 2481
rect 29 2447 45 2481
rect 1213 2447 1229 2481
rect 1287 2447 1303 2481
rect 2471 2447 2487 2481
rect 2545 2447 2561 2481
rect 3729 2447 3745 2481
rect 3803 2447 3819 2481
rect 4987 2447 5003 2481
rect 5061 2447 5077 2481
rect 6245 2447 6261 2481
rect 6319 2447 6335 2481
rect 7503 2447 7519 2481
rect 7577 2447 7593 2481
rect 8761 2447 8777 2481
rect 8835 2447 8851 2481
rect 10019 2447 10035 2481
rect -10081 2388 -10047 2404
rect -10081 -2404 -10047 -2388
rect -8823 2388 -8789 2404
rect -8823 -2404 -8789 -2388
rect -7565 2388 -7531 2404
rect -7565 -2404 -7531 -2388
rect -6307 2388 -6273 2404
rect -6307 -2404 -6273 -2388
rect -5049 2388 -5015 2404
rect -5049 -2404 -5015 -2388
rect -3791 2388 -3757 2404
rect -3791 -2404 -3757 -2388
rect -2533 2388 -2499 2404
rect -2533 -2404 -2499 -2388
rect -1275 2388 -1241 2404
rect -1275 -2404 -1241 -2388
rect -17 2388 17 2404
rect -17 -2404 17 -2388
rect 1241 2388 1275 2404
rect 1241 -2404 1275 -2388
rect 2499 2388 2533 2404
rect 2499 -2404 2533 -2388
rect 3757 2388 3791 2404
rect 3757 -2404 3791 -2388
rect 5015 2388 5049 2404
rect 5015 -2404 5049 -2388
rect 6273 2388 6307 2404
rect 6273 -2404 6307 -2388
rect 7531 2388 7565 2404
rect 7531 -2404 7565 -2388
rect 8789 2388 8823 2404
rect 8789 -2404 8823 -2388
rect 10047 2388 10081 2404
rect 10047 -2404 10081 -2388
rect -10035 -2481 -10019 -2447
rect -8851 -2481 -8835 -2447
rect -8777 -2481 -8761 -2447
rect -7593 -2481 -7577 -2447
rect -7519 -2481 -7503 -2447
rect -6335 -2481 -6319 -2447
rect -6261 -2481 -6245 -2447
rect -5077 -2481 -5061 -2447
rect -5003 -2481 -4987 -2447
rect -3819 -2481 -3803 -2447
rect -3745 -2481 -3729 -2447
rect -2561 -2481 -2545 -2447
rect -2487 -2481 -2471 -2447
rect -1303 -2481 -1287 -2447
rect -1229 -2481 -1213 -2447
rect -45 -2481 -29 -2447
rect 29 -2481 45 -2447
rect 1213 -2481 1229 -2447
rect 1287 -2481 1303 -2447
rect 2471 -2481 2487 -2447
rect 2545 -2481 2561 -2447
rect 3729 -2481 3745 -2447
rect 3803 -2481 3819 -2447
rect 4987 -2481 5003 -2447
rect 5061 -2481 5077 -2447
rect 6245 -2481 6261 -2447
rect 6319 -2481 6335 -2447
rect 7503 -2481 7519 -2447
rect 7577 -2481 7593 -2447
rect 8761 -2481 8777 -2447
rect 8835 -2481 8851 -2447
rect 10019 -2481 10035 -2447
rect -10215 -2585 -10181 -2523
rect 10181 -2585 10215 -2523
rect -10215 -2619 -10119 -2585
rect 10119 -2619 10215 -2585
<< viali >>
rect -10019 2447 -8851 2481
rect -8761 2447 -7593 2481
rect -7503 2447 -6335 2481
rect -6245 2447 -5077 2481
rect -4987 2447 -3819 2481
rect -3729 2447 -2561 2481
rect -2471 2447 -1303 2481
rect -1213 2447 -45 2481
rect 45 2447 1213 2481
rect 1303 2447 2471 2481
rect 2561 2447 3729 2481
rect 3819 2447 4987 2481
rect 5077 2447 6245 2481
rect 6335 2447 7503 2481
rect 7593 2447 8761 2481
rect 8851 2447 10019 2481
rect -10081 -2388 -10047 2388
rect -8823 -2388 -8789 2388
rect -7565 -2388 -7531 2388
rect -6307 -2388 -6273 2388
rect -5049 -2388 -5015 2388
rect -3791 -2388 -3757 2388
rect -2533 -2388 -2499 2388
rect -1275 -2388 -1241 2388
rect -17 -2388 17 2388
rect 1241 -2388 1275 2388
rect 2499 -2388 2533 2388
rect 3757 -2388 3791 2388
rect 5015 -2388 5049 2388
rect 6273 -2388 6307 2388
rect 7531 -2388 7565 2388
rect 8789 -2388 8823 2388
rect 10047 -2388 10081 2388
rect -10019 -2481 -8851 -2447
rect -8761 -2481 -7593 -2447
rect -7503 -2481 -6335 -2447
rect -6245 -2481 -5077 -2447
rect -4987 -2481 -3819 -2447
rect -3729 -2481 -2561 -2447
rect -2471 -2481 -1303 -2447
rect -1213 -2481 -45 -2447
rect 45 -2481 1213 -2447
rect 1303 -2481 2471 -2447
rect 2561 -2481 3729 -2447
rect 3819 -2481 4987 -2447
rect 5077 -2481 6245 -2447
rect 6335 -2481 7503 -2447
rect 7593 -2481 8761 -2447
rect 8851 -2481 10019 -2447
<< metal1 >>
rect -10031 2481 -8839 2487
rect -10031 2447 -10019 2481
rect -8851 2447 -8839 2481
rect -10031 2441 -8839 2447
rect -8773 2481 -7581 2487
rect -8773 2447 -8761 2481
rect -7593 2447 -7581 2481
rect -8773 2441 -7581 2447
rect -7515 2481 -6323 2487
rect -7515 2447 -7503 2481
rect -6335 2447 -6323 2481
rect -7515 2441 -6323 2447
rect -6257 2481 -5065 2487
rect -6257 2447 -6245 2481
rect -5077 2447 -5065 2481
rect -6257 2441 -5065 2447
rect -4999 2481 -3807 2487
rect -4999 2447 -4987 2481
rect -3819 2447 -3807 2481
rect -4999 2441 -3807 2447
rect -3741 2481 -2549 2487
rect -3741 2447 -3729 2481
rect -2561 2447 -2549 2481
rect -3741 2441 -2549 2447
rect -2483 2481 -1291 2487
rect -2483 2447 -2471 2481
rect -1303 2447 -1291 2481
rect -2483 2441 -1291 2447
rect -1225 2481 -33 2487
rect -1225 2447 -1213 2481
rect -45 2447 -33 2481
rect -1225 2441 -33 2447
rect 33 2481 1225 2487
rect 33 2447 45 2481
rect 1213 2447 1225 2481
rect 33 2441 1225 2447
rect 1291 2481 2483 2487
rect 1291 2447 1303 2481
rect 2471 2447 2483 2481
rect 1291 2441 2483 2447
rect 2549 2481 3741 2487
rect 2549 2447 2561 2481
rect 3729 2447 3741 2481
rect 2549 2441 3741 2447
rect 3807 2481 4999 2487
rect 3807 2447 3819 2481
rect 4987 2447 4999 2481
rect 3807 2441 4999 2447
rect 5065 2481 6257 2487
rect 5065 2447 5077 2481
rect 6245 2447 6257 2481
rect 5065 2441 6257 2447
rect 6323 2481 7515 2487
rect 6323 2447 6335 2481
rect 7503 2447 7515 2481
rect 6323 2441 7515 2447
rect 7581 2481 8773 2487
rect 7581 2447 7593 2481
rect 8761 2447 8773 2481
rect 7581 2441 8773 2447
rect 8839 2481 10031 2487
rect 8839 2447 8851 2481
rect 10019 2447 10031 2481
rect 8839 2441 10031 2447
rect -10087 2388 -10041 2400
rect -10087 -2388 -10081 2388
rect -10047 -2388 -10041 2388
rect -10087 -2400 -10041 -2388
rect -8829 2388 -8783 2400
rect -8829 -2388 -8823 2388
rect -8789 -2388 -8783 2388
rect -8829 -2400 -8783 -2388
rect -7571 2388 -7525 2400
rect -7571 -2388 -7565 2388
rect -7531 -2388 -7525 2388
rect -7571 -2400 -7525 -2388
rect -6313 2388 -6267 2400
rect -6313 -2388 -6307 2388
rect -6273 -2388 -6267 2388
rect -6313 -2400 -6267 -2388
rect -5055 2388 -5009 2400
rect -5055 -2388 -5049 2388
rect -5015 -2388 -5009 2388
rect -5055 -2400 -5009 -2388
rect -3797 2388 -3751 2400
rect -3797 -2388 -3791 2388
rect -3757 -2388 -3751 2388
rect -3797 -2400 -3751 -2388
rect -2539 2388 -2493 2400
rect -2539 -2388 -2533 2388
rect -2499 -2388 -2493 2388
rect -2539 -2400 -2493 -2388
rect -1281 2388 -1235 2400
rect -1281 -2388 -1275 2388
rect -1241 -2388 -1235 2388
rect -1281 -2400 -1235 -2388
rect -23 2388 23 2400
rect -23 -2388 -17 2388
rect 17 -2388 23 2388
rect -23 -2400 23 -2388
rect 1235 2388 1281 2400
rect 1235 -2388 1241 2388
rect 1275 -2388 1281 2388
rect 1235 -2400 1281 -2388
rect 2493 2388 2539 2400
rect 2493 -2388 2499 2388
rect 2533 -2388 2539 2388
rect 2493 -2400 2539 -2388
rect 3751 2388 3797 2400
rect 3751 -2388 3757 2388
rect 3791 -2388 3797 2388
rect 3751 -2400 3797 -2388
rect 5009 2388 5055 2400
rect 5009 -2388 5015 2388
rect 5049 -2388 5055 2388
rect 5009 -2400 5055 -2388
rect 6267 2388 6313 2400
rect 6267 -2388 6273 2388
rect 6307 -2388 6313 2388
rect 6267 -2400 6313 -2388
rect 7525 2388 7571 2400
rect 7525 -2388 7531 2388
rect 7565 -2388 7571 2388
rect 7525 -2400 7571 -2388
rect 8783 2388 8829 2400
rect 8783 -2388 8789 2388
rect 8823 -2388 8829 2388
rect 8783 -2400 8829 -2388
rect 10041 2388 10087 2400
rect 10041 -2388 10047 2388
rect 10081 -2388 10087 2388
rect 10041 -2400 10087 -2388
rect -10031 -2447 -8839 -2441
rect -10031 -2481 -10019 -2447
rect -8851 -2481 -8839 -2447
rect -10031 -2487 -8839 -2481
rect -8773 -2447 -7581 -2441
rect -8773 -2481 -8761 -2447
rect -7593 -2481 -7581 -2447
rect -8773 -2487 -7581 -2481
rect -7515 -2447 -6323 -2441
rect -7515 -2481 -7503 -2447
rect -6335 -2481 -6323 -2447
rect -7515 -2487 -6323 -2481
rect -6257 -2447 -5065 -2441
rect -6257 -2481 -6245 -2447
rect -5077 -2481 -5065 -2447
rect -6257 -2487 -5065 -2481
rect -4999 -2447 -3807 -2441
rect -4999 -2481 -4987 -2447
rect -3819 -2481 -3807 -2447
rect -4999 -2487 -3807 -2481
rect -3741 -2447 -2549 -2441
rect -3741 -2481 -3729 -2447
rect -2561 -2481 -2549 -2447
rect -3741 -2487 -2549 -2481
rect -2483 -2447 -1291 -2441
rect -2483 -2481 -2471 -2447
rect -1303 -2481 -1291 -2447
rect -2483 -2487 -1291 -2481
rect -1225 -2447 -33 -2441
rect -1225 -2481 -1213 -2447
rect -45 -2481 -33 -2447
rect -1225 -2487 -33 -2481
rect 33 -2447 1225 -2441
rect 33 -2481 45 -2447
rect 1213 -2481 1225 -2447
rect 33 -2487 1225 -2481
rect 1291 -2447 2483 -2441
rect 1291 -2481 1303 -2447
rect 2471 -2481 2483 -2447
rect 1291 -2487 2483 -2481
rect 2549 -2447 3741 -2441
rect 2549 -2481 2561 -2447
rect 3729 -2481 3741 -2447
rect 2549 -2487 3741 -2481
rect 3807 -2447 4999 -2441
rect 3807 -2481 3819 -2447
rect 4987 -2481 4999 -2447
rect 3807 -2487 4999 -2481
rect 5065 -2447 6257 -2441
rect 5065 -2481 5077 -2447
rect 6245 -2481 6257 -2447
rect 5065 -2487 6257 -2481
rect 6323 -2447 7515 -2441
rect 6323 -2481 6335 -2447
rect 7503 -2481 7515 -2447
rect 6323 -2487 7515 -2481
rect 7581 -2447 8773 -2441
rect 7581 -2481 7593 -2447
rect 8761 -2481 8773 -2447
rect 7581 -2487 8773 -2481
rect 8839 -2447 10031 -2441
rect 8839 -2481 8851 -2447
rect 10019 -2481 10031 -2447
rect 8839 -2487 10031 -2481
<< properties >>
string FIXED_BBOX -10198 -2602 10198 2602
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 24.0 l 6.0 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
