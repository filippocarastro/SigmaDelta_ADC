magic
tech sky130B
magscale 1 2
timestamp 1667224913
<< pwell >>
rect -796 -2579 796 2579
<< nmos >>
rect -600 -2369 600 2431
<< ndiff >>
rect -658 1941 -600 2431
rect -658 -1879 -646 1941
rect -612 -1879 -600 1941
rect -658 -2369 -600 -1879
rect 600 1941 658 2431
rect 600 -1879 612 1941
rect 646 -1879 658 1941
rect 600 -2369 658 -1879
<< ndiffc >>
rect -646 -1879 -612 1941
rect 612 -1879 646 1941
<< psubdiff >>
rect -760 2509 -531 2543
rect 531 2509 760 2543
rect -760 1958 -726 2509
rect -760 -2509 -726 -1958
rect 726 1958 760 2509
rect 726 -2509 760 -1958
rect -760 -2543 -531 -2509
rect 531 -2543 760 -2509
<< psubdiffcont >>
rect -531 2509 531 2543
rect -760 -1958 -726 1958
rect 726 -1958 760 1958
rect -531 -2543 531 -2509
<< poly >>
rect -600 2431 600 2457
rect -600 -2407 600 -2369
rect -600 -2424 -526 -2407
rect -542 -2441 -526 -2424
rect 526 -2424 600 -2407
rect 526 -2441 542 -2424
rect -542 -2457 542 -2441
<< polycont >>
rect -526 -2441 526 -2407
<< locali >>
rect -760 2509 -531 2543
rect 531 2509 760 2543
rect -760 1958 -726 2509
rect 726 1958 760 2509
rect -646 1941 -612 1957
rect -646 -1895 -612 -1879
rect 612 1941 646 1957
rect 612 -1895 646 -1879
rect -760 -2509 -726 -1958
rect -542 -2441 -526 -2407
rect 526 -2441 542 -2407
rect 726 -2509 760 -1958
rect -760 -2543 -531 -2509
rect 531 -2543 760 -2509
<< viali >>
rect -646 -1879 -612 1941
rect 612 -1879 646 1941
rect -526 -2441 526 -2407
<< metal1 >>
rect -652 1941 -606 1953
rect -652 -1879 -646 1941
rect -612 -1879 -606 1941
rect -652 -1891 -606 -1879
rect 606 1941 652 1953
rect 606 -1879 612 1941
rect 646 -1879 652 1941
rect 606 -1891 652 -1879
rect -538 -2407 538 -2401
rect -538 -2441 -526 -2407
rect 526 -2441 538 -2407
rect -538 -2447 538 -2441
<< properties >>
string FIXED_BBOX -743 -2526 743 2526
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 24 l 6 m 1 nf 1 diffcov 80 polycov 90 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 80 rlcov 80 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 80 viadrn 80 viagate 90 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
