magic
tech sky130B
magscale 1 2
timestamp 1667934731
<< nwell >>
rect -4003 -3462 4003 3462
<< mvpmos >>
rect -3745 -3236 -2545 3164
rect -2487 -3236 -1287 3164
rect -1229 -3236 -29 3164
rect 29 -3236 1229 3164
rect 1287 -3236 2487 3164
rect 2545 -3236 3745 3164
<< mvpdiff >>
rect -3803 2514 -3745 3164
rect -3803 -2586 -3791 2514
rect -3757 -2586 -3745 2514
rect -3803 -3236 -3745 -2586
rect -2545 2514 -2487 3164
rect -2545 -2586 -2533 2514
rect -2499 -2586 -2487 2514
rect -2545 -3236 -2487 -2586
rect -1287 2514 -1229 3164
rect -1287 -2586 -1275 2514
rect -1241 -2586 -1229 2514
rect -1287 -3236 -1229 -2586
rect -29 2514 29 3164
rect -29 -2586 -17 2514
rect 17 -2586 29 2514
rect -29 -3236 29 -2586
rect 1229 2514 1287 3164
rect 1229 -2586 1241 2514
rect 1275 -2586 1287 2514
rect 1229 -3236 1287 -2586
rect 2487 2514 2545 3164
rect 2487 -2586 2499 2514
rect 2533 -2586 2545 2514
rect 2487 -3236 2545 -2586
rect 3745 2514 3803 3164
rect 3745 -2586 3757 2514
rect 3791 -2586 3803 2514
rect 3745 -3236 3803 -2586
<< mvpdiffc >>
rect -3791 -2586 -3757 2514
rect -2533 -2586 -2499 2514
rect -1275 -2586 -1241 2514
rect -17 -2586 17 2514
rect 1241 -2586 1275 2514
rect 2499 -2586 2533 2514
rect 3757 -2586 3791 2514
<< mvnsubdiff >>
rect -3937 3338 3937 3396
rect -3937 -3338 -3879 3338
rect 3879 -3338 3937 3338
rect -3937 -3396 3937 -3338
<< poly >>
rect -3687 3245 -2603 3261
rect -3687 3228 -3671 3245
rect -3745 3211 -3671 3228
rect -2619 3228 -2603 3245
rect -2429 3245 -1345 3261
rect -2429 3228 -2413 3245
rect -2619 3211 -2545 3228
rect -3745 3164 -2545 3211
rect -2487 3211 -2413 3228
rect -1361 3228 -1345 3245
rect -1171 3245 -87 3261
rect -1171 3228 -1155 3245
rect -1361 3211 -1287 3228
rect -2487 3164 -1287 3211
rect -1229 3211 -1155 3228
rect -103 3228 -87 3245
rect 87 3245 1171 3261
rect 87 3228 103 3245
rect -103 3211 -29 3228
rect -1229 3164 -29 3211
rect 29 3211 103 3228
rect 1155 3228 1171 3245
rect 1345 3245 2429 3261
rect 1345 3228 1361 3245
rect 1155 3211 1229 3228
rect 29 3164 1229 3211
rect 1287 3211 1361 3228
rect 2413 3228 2429 3245
rect 2603 3245 3687 3261
rect 2603 3228 2619 3245
rect 2413 3211 2487 3228
rect 1287 3164 2487 3211
rect 2545 3211 2619 3228
rect 3671 3228 3687 3245
rect 3671 3211 3745 3228
rect 2545 3164 3745 3211
rect -3745 -3262 -2545 -3236
rect -2487 -3262 -1287 -3236
rect -1229 -3262 -29 -3236
rect 29 -3262 1229 -3236
rect 1287 -3262 2487 -3236
rect 2545 -3262 3745 -3236
<< polycont >>
rect -3671 3211 -2619 3245
rect -2413 3211 -1361 3245
rect -1155 3211 -103 3245
rect 103 3211 1155 3245
rect 1361 3211 2413 3245
rect 2619 3211 3671 3245
<< locali >>
rect -3687 3211 -3671 3245
rect -2619 3211 -2603 3245
rect -2429 3211 -2413 3245
rect -1361 3211 -1345 3245
rect -1171 3211 -1155 3245
rect -103 3211 -87 3245
rect 87 3211 103 3245
rect 1155 3211 1171 3245
rect 1345 3211 1361 3245
rect 2413 3211 2429 3245
rect 2603 3211 2619 3245
rect 3671 3211 3687 3245
rect -3791 2514 -3757 2530
rect -3791 -2602 -3757 -2586
rect -2533 2514 -2499 2530
rect -2533 -2602 -2499 -2586
rect -1275 2514 -1241 2530
rect -1275 -2602 -1241 -2586
rect -17 2514 17 2530
rect -17 -2602 17 -2586
rect 1241 2514 1275 2530
rect 1241 -2602 1275 -2586
rect 2499 2514 2533 2530
rect 2499 -2602 2533 -2586
rect 3757 2514 3791 2530
rect 3757 -2602 3791 -2586
<< viali >>
rect -3671 3211 -2619 3245
rect -2413 3211 -1361 3245
rect -1155 3211 -103 3245
rect 103 3211 1155 3245
rect 1361 3211 2413 3245
rect 2619 3211 3671 3245
rect -3791 -2586 -3757 2514
rect -2533 -2586 -2499 2514
rect -1275 -2586 -1241 2514
rect -17 -2586 17 2514
rect 1241 -2586 1275 2514
rect 2499 -2586 2533 2514
rect 3757 -2586 3791 2514
<< metal1 >>
rect -3683 3245 -2607 3251
rect -3683 3211 -3671 3245
rect -2619 3211 -2607 3245
rect -3683 3205 -2607 3211
rect -2425 3245 -1349 3251
rect -2425 3211 -2413 3245
rect -1361 3211 -1349 3245
rect -2425 3205 -1349 3211
rect -1167 3245 -91 3251
rect -1167 3211 -1155 3245
rect -103 3211 -91 3245
rect -1167 3205 -91 3211
rect 91 3245 1167 3251
rect 91 3211 103 3245
rect 1155 3211 1167 3245
rect 91 3205 1167 3211
rect 1349 3245 2425 3251
rect 1349 3211 1361 3245
rect 2413 3211 2425 3245
rect 1349 3205 2425 3211
rect 2607 3245 3683 3251
rect 2607 3211 2619 3245
rect 3671 3211 3683 3245
rect 2607 3205 3683 3211
rect -3797 2514 -3751 2526
rect -3797 -2586 -3791 2514
rect -3757 -2586 -3751 2514
rect -3797 -2598 -3751 -2586
rect -2539 2514 -2493 2526
rect -2539 -2586 -2533 2514
rect -2499 -2586 -2493 2514
rect -2539 -2598 -2493 -2586
rect -1281 2514 -1235 2526
rect -1281 -2586 -1275 2514
rect -1241 -2586 -1235 2514
rect -1281 -2598 -1235 -2586
rect -23 2514 23 2526
rect -23 -2586 -17 2514
rect 17 -2586 23 2514
rect -23 -2598 23 -2586
rect 1235 2514 1281 2526
rect 1235 -2586 1241 2514
rect 1275 -2586 1281 2514
rect 1235 -2598 1281 -2586
rect 2493 2514 2539 2526
rect 2493 -2586 2499 2514
rect 2533 -2586 2539 2514
rect 2493 -2598 2539 -2586
rect 3751 2514 3797 2526
rect 3751 -2586 3757 2514
rect 3791 -2586 3797 2514
rect 3751 -2598 3797 -2586
<< properties >>
string FIXED_BBOX -3908 -3367 3908 3367
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 6.0 m 1 nf 6 diffcov 80 polycov 90 guard 1 glc 0 grc 0 gtc 0 gbc 0 tbcov 80 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 80 viadrn 80 viagate 90 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
