magic
tech sky130B
magscale 1 2
timestamp 1667069824
<< nwell >>
rect -10293 -2662 10293 2662
<< mvpmos >>
rect -10035 -2436 -8835 2364
rect -8777 -2436 -7577 2364
rect -7519 -2436 -6319 2364
rect -6261 -2436 -5061 2364
rect -5003 -2436 -3803 2364
rect -3745 -2436 -2545 2364
rect -2487 -2436 -1287 2364
rect -1229 -2436 -29 2364
rect 29 -2436 1229 2364
rect 1287 -2436 2487 2364
rect 2545 -2436 3745 2364
rect 3803 -2436 5003 2364
rect 5061 -2436 6261 2364
rect 6319 -2436 7519 2364
rect 7577 -2436 8777 2364
rect 8835 -2436 10035 2364
<< mvpdiff >>
rect -10093 2352 -10035 2364
rect -10093 -2424 -10081 2352
rect -10047 -2424 -10035 2352
rect -10093 -2436 -10035 -2424
rect -8835 2352 -8777 2364
rect -8835 -2424 -8823 2352
rect -8789 -2424 -8777 2352
rect -8835 -2436 -8777 -2424
rect -7577 2352 -7519 2364
rect -7577 -2424 -7565 2352
rect -7531 -2424 -7519 2352
rect -7577 -2436 -7519 -2424
rect -6319 2352 -6261 2364
rect -6319 -2424 -6307 2352
rect -6273 -2424 -6261 2352
rect -6319 -2436 -6261 -2424
rect -5061 2352 -5003 2364
rect -5061 -2424 -5049 2352
rect -5015 -2424 -5003 2352
rect -5061 -2436 -5003 -2424
rect -3803 2352 -3745 2364
rect -3803 -2424 -3791 2352
rect -3757 -2424 -3745 2352
rect -3803 -2436 -3745 -2424
rect -2545 2352 -2487 2364
rect -2545 -2424 -2533 2352
rect -2499 -2424 -2487 2352
rect -2545 -2436 -2487 -2424
rect -1287 2352 -1229 2364
rect -1287 -2424 -1275 2352
rect -1241 -2424 -1229 2352
rect -1287 -2436 -1229 -2424
rect -29 2352 29 2364
rect -29 -2424 -17 2352
rect 17 -2424 29 2352
rect -29 -2436 29 -2424
rect 1229 2352 1287 2364
rect 1229 -2424 1241 2352
rect 1275 -2424 1287 2352
rect 1229 -2436 1287 -2424
rect 2487 2352 2545 2364
rect 2487 -2424 2499 2352
rect 2533 -2424 2545 2352
rect 2487 -2436 2545 -2424
rect 3745 2352 3803 2364
rect 3745 -2424 3757 2352
rect 3791 -2424 3803 2352
rect 3745 -2436 3803 -2424
rect 5003 2352 5061 2364
rect 5003 -2424 5015 2352
rect 5049 -2424 5061 2352
rect 5003 -2436 5061 -2424
rect 6261 2352 6319 2364
rect 6261 -2424 6273 2352
rect 6307 -2424 6319 2352
rect 6261 -2436 6319 -2424
rect 7519 2352 7577 2364
rect 7519 -2424 7531 2352
rect 7565 -2424 7577 2352
rect 7519 -2436 7577 -2424
rect 8777 2352 8835 2364
rect 8777 -2424 8789 2352
rect 8823 -2424 8835 2352
rect 8777 -2436 8835 -2424
rect 10035 2352 10093 2364
rect 10035 -2424 10047 2352
rect 10081 -2424 10093 2352
rect 10035 -2436 10093 -2424
<< mvpdiffc >>
rect -10081 -2424 -10047 2352
rect -8823 -2424 -8789 2352
rect -7565 -2424 -7531 2352
rect -6307 -2424 -6273 2352
rect -5049 -2424 -5015 2352
rect -3791 -2424 -3757 2352
rect -2533 -2424 -2499 2352
rect -1275 -2424 -1241 2352
rect -17 -2424 17 2352
rect 1241 -2424 1275 2352
rect 2499 -2424 2533 2352
rect 3757 -2424 3791 2352
rect 5015 -2424 5049 2352
rect 6273 -2424 6307 2352
rect 7531 -2424 7565 2352
rect 8789 -2424 8823 2352
rect 10047 -2424 10081 2352
<< mvnsubdiff >>
rect -10227 2584 10227 2596
rect -10227 2550 -10119 2584
rect 10119 2550 10227 2584
rect -10227 2538 10227 2550
rect -10227 2488 -10169 2538
rect -10227 -2488 -10215 2488
rect -10181 -2488 -10169 2488
rect 10169 2488 10227 2538
rect -10227 -2538 -10169 -2488
rect 10169 -2488 10181 2488
rect 10215 -2488 10227 2488
rect 10169 -2538 10227 -2488
rect -10227 -2550 10227 -2538
rect -10227 -2584 -10119 -2550
rect 10119 -2584 10227 -2550
rect -10227 -2596 10227 -2584
<< mvnsubdiffcont >>
rect -10119 2550 10119 2584
rect -10215 -2488 -10181 2488
rect 10181 -2488 10215 2488
rect -10119 -2584 10119 -2550
<< poly >>
rect -10035 2445 -8835 2461
rect -10035 2411 -10019 2445
rect -8851 2411 -8835 2445
rect -10035 2364 -8835 2411
rect -8777 2445 -7577 2461
rect -8777 2411 -8761 2445
rect -7593 2411 -7577 2445
rect -8777 2364 -7577 2411
rect -7519 2445 -6319 2461
rect -7519 2411 -7503 2445
rect -6335 2411 -6319 2445
rect -7519 2364 -6319 2411
rect -6261 2445 -5061 2461
rect -6261 2411 -6245 2445
rect -5077 2411 -5061 2445
rect -6261 2364 -5061 2411
rect -5003 2445 -3803 2461
rect -5003 2411 -4987 2445
rect -3819 2411 -3803 2445
rect -5003 2364 -3803 2411
rect -3745 2445 -2545 2461
rect -3745 2411 -3729 2445
rect -2561 2411 -2545 2445
rect -3745 2364 -2545 2411
rect -2487 2445 -1287 2461
rect -2487 2411 -2471 2445
rect -1303 2411 -1287 2445
rect -2487 2364 -1287 2411
rect -1229 2445 -29 2461
rect -1229 2411 -1213 2445
rect -45 2411 -29 2445
rect -1229 2364 -29 2411
rect 29 2445 1229 2461
rect 29 2411 45 2445
rect 1213 2411 1229 2445
rect 29 2364 1229 2411
rect 1287 2445 2487 2461
rect 1287 2411 1303 2445
rect 2471 2411 2487 2445
rect 1287 2364 2487 2411
rect 2545 2445 3745 2461
rect 2545 2411 2561 2445
rect 3729 2411 3745 2445
rect 2545 2364 3745 2411
rect 3803 2445 5003 2461
rect 3803 2411 3819 2445
rect 4987 2411 5003 2445
rect 3803 2364 5003 2411
rect 5061 2445 6261 2461
rect 5061 2411 5077 2445
rect 6245 2411 6261 2445
rect 5061 2364 6261 2411
rect 6319 2445 7519 2461
rect 6319 2411 6335 2445
rect 7503 2411 7519 2445
rect 6319 2364 7519 2411
rect 7577 2445 8777 2461
rect 7577 2411 7593 2445
rect 8761 2411 8777 2445
rect 7577 2364 8777 2411
rect 8835 2445 10035 2461
rect 8835 2411 8851 2445
rect 10019 2411 10035 2445
rect 8835 2364 10035 2411
rect -10035 -2462 -8835 -2436
rect -8777 -2462 -7577 -2436
rect -7519 -2462 -6319 -2436
rect -6261 -2462 -5061 -2436
rect -5003 -2462 -3803 -2436
rect -3745 -2462 -2545 -2436
rect -2487 -2462 -1287 -2436
rect -1229 -2462 -29 -2436
rect 29 -2462 1229 -2436
rect 1287 -2462 2487 -2436
rect 2545 -2462 3745 -2436
rect 3803 -2462 5003 -2436
rect 5061 -2462 6261 -2436
rect 6319 -2462 7519 -2436
rect 7577 -2462 8777 -2436
rect 8835 -2462 10035 -2436
<< polycont >>
rect -10019 2411 -8851 2445
rect -8761 2411 -7593 2445
rect -7503 2411 -6335 2445
rect -6245 2411 -5077 2445
rect -4987 2411 -3819 2445
rect -3729 2411 -2561 2445
rect -2471 2411 -1303 2445
rect -1213 2411 -45 2445
rect 45 2411 1213 2445
rect 1303 2411 2471 2445
rect 2561 2411 3729 2445
rect 3819 2411 4987 2445
rect 5077 2411 6245 2445
rect 6335 2411 7503 2445
rect 7593 2411 8761 2445
rect 8851 2411 10019 2445
<< locali >>
rect -10215 2550 -10119 2584
rect 10119 2550 10215 2584
rect -10215 2488 -10181 2550
rect 10181 2488 10215 2550
rect -10035 2411 -10019 2445
rect -8851 2411 -8835 2445
rect -8777 2411 -8761 2445
rect -7593 2411 -7577 2445
rect -7519 2411 -7503 2445
rect -6335 2411 -6319 2445
rect -6261 2411 -6245 2445
rect -5077 2411 -5061 2445
rect -5003 2411 -4987 2445
rect -3819 2411 -3803 2445
rect -3745 2411 -3729 2445
rect -2561 2411 -2545 2445
rect -2487 2411 -2471 2445
rect -1303 2411 -1287 2445
rect -1229 2411 -1213 2445
rect -45 2411 -29 2445
rect 29 2411 45 2445
rect 1213 2411 1229 2445
rect 1287 2411 1303 2445
rect 2471 2411 2487 2445
rect 2545 2411 2561 2445
rect 3729 2411 3745 2445
rect 3803 2411 3819 2445
rect 4987 2411 5003 2445
rect 5061 2411 5077 2445
rect 6245 2411 6261 2445
rect 6319 2411 6335 2445
rect 7503 2411 7519 2445
rect 7577 2411 7593 2445
rect 8761 2411 8777 2445
rect 8835 2411 8851 2445
rect 10019 2411 10035 2445
rect -10081 2352 -10047 2368
rect -10081 -2440 -10047 -2424
rect -8823 2352 -8789 2368
rect -8823 -2440 -8789 -2424
rect -7565 2352 -7531 2368
rect -7565 -2440 -7531 -2424
rect -6307 2352 -6273 2368
rect -6307 -2440 -6273 -2424
rect -5049 2352 -5015 2368
rect -5049 -2440 -5015 -2424
rect -3791 2352 -3757 2368
rect -3791 -2440 -3757 -2424
rect -2533 2352 -2499 2368
rect -2533 -2440 -2499 -2424
rect -1275 2352 -1241 2368
rect -1275 -2440 -1241 -2424
rect -17 2352 17 2368
rect -17 -2440 17 -2424
rect 1241 2352 1275 2368
rect 1241 -2440 1275 -2424
rect 2499 2352 2533 2368
rect 2499 -2440 2533 -2424
rect 3757 2352 3791 2368
rect 3757 -2440 3791 -2424
rect 5015 2352 5049 2368
rect 5015 -2440 5049 -2424
rect 6273 2352 6307 2368
rect 6273 -2440 6307 -2424
rect 7531 2352 7565 2368
rect 7531 -2440 7565 -2424
rect 8789 2352 8823 2368
rect 8789 -2440 8823 -2424
rect 10047 2352 10081 2368
rect 10047 -2440 10081 -2424
rect -10215 -2550 -10181 -2488
rect 10181 -2550 10215 -2488
rect -10215 -2584 -10119 -2550
rect 10119 -2584 10215 -2550
<< viali >>
rect -10019 2411 -8851 2445
rect -8761 2411 -7593 2445
rect -7503 2411 -6335 2445
rect -6245 2411 -5077 2445
rect -4987 2411 -3819 2445
rect -3729 2411 -2561 2445
rect -2471 2411 -1303 2445
rect -1213 2411 -45 2445
rect 45 2411 1213 2445
rect 1303 2411 2471 2445
rect 2561 2411 3729 2445
rect 3819 2411 4987 2445
rect 5077 2411 6245 2445
rect 6335 2411 7503 2445
rect 7593 2411 8761 2445
rect 8851 2411 10019 2445
rect -10081 -2424 -10047 2352
rect -8823 -2424 -8789 2352
rect -7565 -2424 -7531 2352
rect -6307 -2424 -6273 2352
rect -5049 -2424 -5015 2352
rect -3791 -2424 -3757 2352
rect -2533 -2424 -2499 2352
rect -1275 -2424 -1241 2352
rect -17 -2424 17 2352
rect 1241 -2424 1275 2352
rect 2499 -2424 2533 2352
rect 3757 -2424 3791 2352
rect 5015 -2424 5049 2352
rect 6273 -2424 6307 2352
rect 7531 -2424 7565 2352
rect 8789 -2424 8823 2352
rect 10047 -2424 10081 2352
<< metal1 >>
rect -10031 2445 -8839 2451
rect -10031 2411 -10019 2445
rect -8851 2411 -8839 2445
rect -10031 2405 -8839 2411
rect -8773 2445 -7581 2451
rect -8773 2411 -8761 2445
rect -7593 2411 -7581 2445
rect -8773 2405 -7581 2411
rect -7515 2445 -6323 2451
rect -7515 2411 -7503 2445
rect -6335 2411 -6323 2445
rect -7515 2405 -6323 2411
rect -6257 2445 -5065 2451
rect -6257 2411 -6245 2445
rect -5077 2411 -5065 2445
rect -6257 2405 -5065 2411
rect -4999 2445 -3807 2451
rect -4999 2411 -4987 2445
rect -3819 2411 -3807 2445
rect -4999 2405 -3807 2411
rect -3741 2445 -2549 2451
rect -3741 2411 -3729 2445
rect -2561 2411 -2549 2445
rect -3741 2405 -2549 2411
rect -2483 2445 -1291 2451
rect -2483 2411 -2471 2445
rect -1303 2411 -1291 2445
rect -2483 2405 -1291 2411
rect -1225 2445 -33 2451
rect -1225 2411 -1213 2445
rect -45 2411 -33 2445
rect -1225 2405 -33 2411
rect 33 2445 1225 2451
rect 33 2411 45 2445
rect 1213 2411 1225 2445
rect 33 2405 1225 2411
rect 1291 2445 2483 2451
rect 1291 2411 1303 2445
rect 2471 2411 2483 2445
rect 1291 2405 2483 2411
rect 2549 2445 3741 2451
rect 2549 2411 2561 2445
rect 3729 2411 3741 2445
rect 2549 2405 3741 2411
rect 3807 2445 4999 2451
rect 3807 2411 3819 2445
rect 4987 2411 4999 2445
rect 3807 2405 4999 2411
rect 5065 2445 6257 2451
rect 5065 2411 5077 2445
rect 6245 2411 6257 2445
rect 5065 2405 6257 2411
rect 6323 2445 7515 2451
rect 6323 2411 6335 2445
rect 7503 2411 7515 2445
rect 6323 2405 7515 2411
rect 7581 2445 8773 2451
rect 7581 2411 7593 2445
rect 8761 2411 8773 2445
rect 7581 2405 8773 2411
rect 8839 2445 10031 2451
rect 8839 2411 8851 2445
rect 10019 2411 10031 2445
rect 8839 2405 10031 2411
rect -10087 2352 -10041 2364
rect -10087 -2424 -10081 2352
rect -10047 -2424 -10041 2352
rect -10087 -2436 -10041 -2424
rect -8829 2352 -8783 2364
rect -8829 -2424 -8823 2352
rect -8789 -2424 -8783 2352
rect -8829 -2436 -8783 -2424
rect -7571 2352 -7525 2364
rect -7571 -2424 -7565 2352
rect -7531 -2424 -7525 2352
rect -7571 -2436 -7525 -2424
rect -6313 2352 -6267 2364
rect -6313 -2424 -6307 2352
rect -6273 -2424 -6267 2352
rect -6313 -2436 -6267 -2424
rect -5055 2352 -5009 2364
rect -5055 -2424 -5049 2352
rect -5015 -2424 -5009 2352
rect -5055 -2436 -5009 -2424
rect -3797 2352 -3751 2364
rect -3797 -2424 -3791 2352
rect -3757 -2424 -3751 2352
rect -3797 -2436 -3751 -2424
rect -2539 2352 -2493 2364
rect -2539 -2424 -2533 2352
rect -2499 -2424 -2493 2352
rect -2539 -2436 -2493 -2424
rect -1281 2352 -1235 2364
rect -1281 -2424 -1275 2352
rect -1241 -2424 -1235 2352
rect -1281 -2436 -1235 -2424
rect -23 2352 23 2364
rect -23 -2424 -17 2352
rect 17 -2424 23 2352
rect -23 -2436 23 -2424
rect 1235 2352 1281 2364
rect 1235 -2424 1241 2352
rect 1275 -2424 1281 2352
rect 1235 -2436 1281 -2424
rect 2493 2352 2539 2364
rect 2493 -2424 2499 2352
rect 2533 -2424 2539 2352
rect 2493 -2436 2539 -2424
rect 3751 2352 3797 2364
rect 3751 -2424 3757 2352
rect 3791 -2424 3797 2352
rect 3751 -2436 3797 -2424
rect 5009 2352 5055 2364
rect 5009 -2424 5015 2352
rect 5049 -2424 5055 2352
rect 5009 -2436 5055 -2424
rect 6267 2352 6313 2364
rect 6267 -2424 6273 2352
rect 6307 -2424 6313 2352
rect 6267 -2436 6313 -2424
rect 7525 2352 7571 2364
rect 7525 -2424 7531 2352
rect 7565 -2424 7571 2352
rect 7525 -2436 7571 -2424
rect 8783 2352 8829 2364
rect 8783 -2424 8789 2352
rect 8823 -2424 8829 2352
rect 8783 -2436 8829 -2424
rect 10041 2352 10087 2364
rect 10041 -2424 10047 2352
rect 10081 -2424 10087 2352
rect 10041 -2436 10087 -2424
<< properties >>
string FIXED_BBOX -10198 -2567 10198 2567
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 24.0 l 6.0 m 1 nf 16 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
