magic
tech sky130B
magscale 1 2
timestamp 1667069824
<< nwell >>
rect -858 -19874 858 19874
<< mvpmos >>
rect -600 13177 600 19577
rect -600 6612 600 13012
rect -600 47 600 6447
rect -600 -6518 600 -118
rect -600 -13083 600 -6683
rect -600 -19648 600 -13248
<< mvpdiff >>
rect -658 19565 -600 19577
rect -658 13189 -646 19565
rect -612 13189 -600 19565
rect -658 13177 -600 13189
rect 600 19565 658 19577
rect 600 13189 612 19565
rect 646 13189 658 19565
rect 600 13177 658 13189
rect -658 13000 -600 13012
rect -658 6624 -646 13000
rect -612 6624 -600 13000
rect -658 6612 -600 6624
rect 600 13000 658 13012
rect 600 6624 612 13000
rect 646 6624 658 13000
rect 600 6612 658 6624
rect -658 6435 -600 6447
rect -658 59 -646 6435
rect -612 59 -600 6435
rect -658 47 -600 59
rect 600 6435 658 6447
rect 600 59 612 6435
rect 646 59 658 6435
rect 600 47 658 59
rect -658 -130 -600 -118
rect -658 -6506 -646 -130
rect -612 -6506 -600 -130
rect -658 -6518 -600 -6506
rect 600 -130 658 -118
rect 600 -6506 612 -130
rect 646 -6506 658 -130
rect 600 -6518 658 -6506
rect -658 -6695 -600 -6683
rect -658 -13071 -646 -6695
rect -612 -13071 -600 -6695
rect -658 -13083 -600 -13071
rect 600 -6695 658 -6683
rect 600 -13071 612 -6695
rect 646 -13071 658 -6695
rect 600 -13083 658 -13071
rect -658 -13260 -600 -13248
rect -658 -19636 -646 -13260
rect -612 -19636 -600 -13260
rect -658 -19648 -600 -19636
rect 600 -13260 658 -13248
rect 600 -19636 612 -13260
rect 646 -19636 658 -13260
rect 600 -19648 658 -19636
<< mvpdiffc >>
rect -646 13189 -612 19565
rect 612 13189 646 19565
rect -646 6624 -612 13000
rect 612 6624 646 13000
rect -646 59 -612 6435
rect 612 59 646 6435
rect -646 -6506 -612 -130
rect 612 -6506 646 -130
rect -646 -13071 -612 -6695
rect 612 -13071 646 -6695
rect -646 -19636 -612 -13260
rect 612 -19636 646 -13260
<< mvnsubdiff >>
rect -792 19796 792 19808
rect -792 19762 -684 19796
rect 684 19762 792 19796
rect -792 19750 792 19762
rect -792 19700 -734 19750
rect -792 -19700 -780 19700
rect -746 -19700 -734 19700
rect 734 19700 792 19750
rect -792 -19750 -734 -19700
rect 734 -19700 746 19700
rect 780 -19700 792 19700
rect 734 -19750 792 -19700
rect -792 -19762 792 -19750
rect -792 -19796 -684 -19762
rect 684 -19796 792 -19762
rect -792 -19808 792 -19796
<< mvnsubdiffcont >>
rect -684 19762 684 19796
rect -780 -19700 -746 19700
rect 746 -19700 780 19700
rect -684 -19796 684 -19762
<< poly >>
rect -600 19658 600 19674
rect -600 19624 -584 19658
rect 584 19624 600 19658
rect -600 19577 600 19624
rect -600 13151 600 13177
rect -600 13093 600 13109
rect -600 13059 -584 13093
rect 584 13059 600 13093
rect -600 13012 600 13059
rect -600 6586 600 6612
rect -600 6528 600 6544
rect -600 6494 -584 6528
rect 584 6494 600 6528
rect -600 6447 600 6494
rect -600 21 600 47
rect -600 -37 600 -21
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -600 -118 600 -71
rect -600 -6544 600 -6518
rect -600 -6602 600 -6586
rect -600 -6636 -584 -6602
rect 584 -6636 600 -6602
rect -600 -6683 600 -6636
rect -600 -13109 600 -13083
rect -600 -13167 600 -13151
rect -600 -13201 -584 -13167
rect 584 -13201 600 -13167
rect -600 -13248 600 -13201
rect -600 -19674 600 -19648
<< polycont >>
rect -584 19624 584 19658
rect -584 13059 584 13093
rect -584 6494 584 6528
rect -584 -71 584 -37
rect -584 -6636 584 -6602
rect -584 -13201 584 -13167
<< locali >>
rect -780 19762 -684 19796
rect 684 19762 780 19796
rect -780 19700 -746 19762
rect 746 19700 780 19762
rect -600 19624 -584 19658
rect 584 19624 600 19658
rect -646 19565 -612 19581
rect -646 13173 -612 13189
rect 612 19565 646 19581
rect 612 13173 646 13189
rect -600 13059 -584 13093
rect 584 13059 600 13093
rect -646 13000 -612 13016
rect -646 6608 -612 6624
rect 612 13000 646 13016
rect 612 6608 646 6624
rect -600 6494 -584 6528
rect 584 6494 600 6528
rect -646 6435 -612 6451
rect -646 43 -612 59
rect 612 6435 646 6451
rect 612 43 646 59
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -646 -130 -612 -114
rect -646 -6522 -612 -6506
rect 612 -130 646 -114
rect 612 -6522 646 -6506
rect -600 -6636 -584 -6602
rect 584 -6636 600 -6602
rect -646 -6695 -612 -6679
rect -646 -13087 -612 -13071
rect 612 -6695 646 -6679
rect 612 -13087 646 -13071
rect -600 -13201 -584 -13167
rect 584 -13201 600 -13167
rect -646 -13260 -612 -13244
rect -646 -19652 -612 -19636
rect 612 -13260 646 -13244
rect 612 -19652 646 -19636
rect -780 -19762 -746 -19700
rect 746 -19762 780 -19700
rect -780 -19796 -684 -19762
rect 684 -19796 780 -19762
<< viali >>
rect -584 19624 584 19658
rect -646 13189 -612 19565
rect 612 13189 646 19565
rect -584 13059 584 13093
rect -646 6624 -612 13000
rect 612 6624 646 13000
rect -584 6494 584 6528
rect -646 59 -612 6435
rect 612 59 646 6435
rect -584 -71 584 -37
rect -646 -6506 -612 -130
rect 612 -6506 646 -130
rect -584 -6636 584 -6602
rect -646 -13071 -612 -6695
rect 612 -13071 646 -6695
rect -584 -13201 584 -13167
rect -646 -19636 -612 -13260
rect 612 -19636 646 -13260
<< metal1 >>
rect -596 19658 596 19664
rect -596 19624 -584 19658
rect 584 19624 596 19658
rect -596 19618 596 19624
rect -652 19565 -606 19577
rect -652 13189 -646 19565
rect -612 13189 -606 19565
rect -652 13177 -606 13189
rect 606 19565 652 19577
rect 606 13189 612 19565
rect 646 13189 652 19565
rect 606 13177 652 13189
rect -596 13093 596 13099
rect -596 13059 -584 13093
rect 584 13059 596 13093
rect -596 13053 596 13059
rect -652 13000 -606 13012
rect -652 6624 -646 13000
rect -612 6624 -606 13000
rect -652 6612 -606 6624
rect 606 13000 652 13012
rect 606 6624 612 13000
rect 646 6624 652 13000
rect 606 6612 652 6624
rect -596 6528 596 6534
rect -596 6494 -584 6528
rect 584 6494 596 6528
rect -596 6488 596 6494
rect -652 6435 -606 6447
rect -652 59 -646 6435
rect -612 59 -606 6435
rect -652 47 -606 59
rect 606 6435 652 6447
rect 606 59 612 6435
rect 646 59 652 6435
rect 606 47 652 59
rect -596 -37 596 -31
rect -596 -71 -584 -37
rect 584 -71 596 -37
rect -596 -77 596 -71
rect -652 -130 -606 -118
rect -652 -6506 -646 -130
rect -612 -6506 -606 -130
rect -652 -6518 -606 -6506
rect 606 -130 652 -118
rect 606 -6506 612 -130
rect 646 -6506 652 -130
rect 606 -6518 652 -6506
rect -596 -6602 596 -6596
rect -596 -6636 -584 -6602
rect 584 -6636 596 -6602
rect -596 -6642 596 -6636
rect -652 -6695 -606 -6683
rect -652 -13071 -646 -6695
rect -612 -13071 -606 -6695
rect -652 -13083 -606 -13071
rect 606 -6695 652 -6683
rect 606 -13071 612 -6695
rect 646 -13071 652 -6695
rect 606 -13083 652 -13071
rect -596 -13167 596 -13161
rect -596 -13201 -584 -13167
rect 584 -13201 596 -13167
rect -596 -13207 596 -13201
rect -652 -13260 -606 -13248
rect -652 -19636 -646 -13260
rect -612 -19636 -606 -13260
rect -652 -19648 -606 -19636
rect 606 -13260 652 -13248
rect 606 -19636 612 -13260
rect 646 -19636 652 -13260
rect 606 -19648 652 -19636
<< properties >>
string FIXED_BBOX -763 -19779 763 19779
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 6.0 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
