magic
tech sky130B
magscale 1 2
timestamp 1667069824
<< nwell >>
rect -4003 -3462 4003 3462
<< mvpmos >>
rect -3745 -3236 -2545 3164
rect -2487 -3236 -1287 3164
rect -1229 -3236 -29 3164
rect 29 -3236 1229 3164
rect 1287 -3236 2487 3164
rect 2545 -3236 3745 3164
<< mvpdiff >>
rect -3803 3152 -3745 3164
rect -3803 -3224 -3791 3152
rect -3757 -3224 -3745 3152
rect -3803 -3236 -3745 -3224
rect -2545 3152 -2487 3164
rect -2545 -3224 -2533 3152
rect -2499 -3224 -2487 3152
rect -2545 -3236 -2487 -3224
rect -1287 3152 -1229 3164
rect -1287 -3224 -1275 3152
rect -1241 -3224 -1229 3152
rect -1287 -3236 -1229 -3224
rect -29 3152 29 3164
rect -29 -3224 -17 3152
rect 17 -3224 29 3152
rect -29 -3236 29 -3224
rect 1229 3152 1287 3164
rect 1229 -3224 1241 3152
rect 1275 -3224 1287 3152
rect 1229 -3236 1287 -3224
rect 2487 3152 2545 3164
rect 2487 -3224 2499 3152
rect 2533 -3224 2545 3152
rect 2487 -3236 2545 -3224
rect 3745 3152 3803 3164
rect 3745 -3224 3757 3152
rect 3791 -3224 3803 3152
rect 3745 -3236 3803 -3224
<< mvpdiffc >>
rect -3791 -3224 -3757 3152
rect -2533 -3224 -2499 3152
rect -1275 -3224 -1241 3152
rect -17 -3224 17 3152
rect 1241 -3224 1275 3152
rect 2499 -3224 2533 3152
rect 3757 -3224 3791 3152
<< mvnsubdiff >>
rect -3937 3384 3937 3396
rect -3937 3350 -3829 3384
rect 3829 3350 3937 3384
rect -3937 3338 3937 3350
rect -3937 3288 -3879 3338
rect -3937 -3288 -3925 3288
rect -3891 -3288 -3879 3288
rect 3879 3288 3937 3338
rect -3937 -3338 -3879 -3288
rect 3879 -3288 3891 3288
rect 3925 -3288 3937 3288
rect 3879 -3338 3937 -3288
rect -3937 -3350 3937 -3338
rect -3937 -3384 -3829 -3350
rect 3829 -3384 3937 -3350
rect -3937 -3396 3937 -3384
<< mvnsubdiffcont >>
rect -3829 3350 3829 3384
rect -3925 -3288 -3891 3288
rect 3891 -3288 3925 3288
rect -3829 -3384 3829 -3350
<< poly >>
rect -3745 3245 -2545 3261
rect -3745 3211 -3729 3245
rect -2561 3211 -2545 3245
rect -3745 3164 -2545 3211
rect -2487 3245 -1287 3261
rect -2487 3211 -2471 3245
rect -1303 3211 -1287 3245
rect -2487 3164 -1287 3211
rect -1229 3245 -29 3261
rect -1229 3211 -1213 3245
rect -45 3211 -29 3245
rect -1229 3164 -29 3211
rect 29 3245 1229 3261
rect 29 3211 45 3245
rect 1213 3211 1229 3245
rect 29 3164 1229 3211
rect 1287 3245 2487 3261
rect 1287 3211 1303 3245
rect 2471 3211 2487 3245
rect 1287 3164 2487 3211
rect 2545 3245 3745 3261
rect 2545 3211 2561 3245
rect 3729 3211 3745 3245
rect 2545 3164 3745 3211
rect -3745 -3262 -2545 -3236
rect -2487 -3262 -1287 -3236
rect -1229 -3262 -29 -3236
rect 29 -3262 1229 -3236
rect 1287 -3262 2487 -3236
rect 2545 -3262 3745 -3236
<< polycont >>
rect -3729 3211 -2561 3245
rect -2471 3211 -1303 3245
rect -1213 3211 -45 3245
rect 45 3211 1213 3245
rect 1303 3211 2471 3245
rect 2561 3211 3729 3245
<< locali >>
rect -3925 3350 -3829 3384
rect 3829 3350 3925 3384
rect -3925 3288 -3891 3350
rect 3891 3288 3925 3350
rect -3745 3211 -3729 3245
rect -2561 3211 -2545 3245
rect -2487 3211 -2471 3245
rect -1303 3211 -1287 3245
rect -1229 3211 -1213 3245
rect -45 3211 -29 3245
rect 29 3211 45 3245
rect 1213 3211 1229 3245
rect 1287 3211 1303 3245
rect 2471 3211 2487 3245
rect 2545 3211 2561 3245
rect 3729 3211 3745 3245
rect -3791 3152 -3757 3168
rect -3791 -3240 -3757 -3224
rect -2533 3152 -2499 3168
rect -2533 -3240 -2499 -3224
rect -1275 3152 -1241 3168
rect -1275 -3240 -1241 -3224
rect -17 3152 17 3168
rect -17 -3240 17 -3224
rect 1241 3152 1275 3168
rect 1241 -3240 1275 -3224
rect 2499 3152 2533 3168
rect 2499 -3240 2533 -3224
rect 3757 3152 3791 3168
rect 3757 -3240 3791 -3224
rect -3925 -3350 -3891 -3288
rect 3891 -3350 3925 -3288
rect -3925 -3384 -3829 -3350
rect 3829 -3384 3925 -3350
<< viali >>
rect -3729 3211 -2561 3245
rect -2471 3211 -1303 3245
rect -1213 3211 -45 3245
rect 45 3211 1213 3245
rect 1303 3211 2471 3245
rect 2561 3211 3729 3245
rect -3791 -3224 -3757 3152
rect -2533 -3224 -2499 3152
rect -1275 -3224 -1241 3152
rect -17 -3224 17 3152
rect 1241 -3224 1275 3152
rect 2499 -3224 2533 3152
rect 3757 -3224 3791 3152
<< metal1 >>
rect -3741 3245 -2549 3251
rect -3741 3211 -3729 3245
rect -2561 3211 -2549 3245
rect -3741 3205 -2549 3211
rect -2483 3245 -1291 3251
rect -2483 3211 -2471 3245
rect -1303 3211 -1291 3245
rect -2483 3205 -1291 3211
rect -1225 3245 -33 3251
rect -1225 3211 -1213 3245
rect -45 3211 -33 3245
rect -1225 3205 -33 3211
rect 33 3245 1225 3251
rect 33 3211 45 3245
rect 1213 3211 1225 3245
rect 33 3205 1225 3211
rect 1291 3245 2483 3251
rect 1291 3211 1303 3245
rect 2471 3211 2483 3245
rect 1291 3205 2483 3211
rect 2549 3245 3741 3251
rect 2549 3211 2561 3245
rect 3729 3211 3741 3245
rect 2549 3205 3741 3211
rect -3797 3152 -3751 3164
rect -3797 -3224 -3791 3152
rect -3757 -3224 -3751 3152
rect -3797 -3236 -3751 -3224
rect -2539 3152 -2493 3164
rect -2539 -3224 -2533 3152
rect -2499 -3224 -2493 3152
rect -2539 -3236 -2493 -3224
rect -1281 3152 -1235 3164
rect -1281 -3224 -1275 3152
rect -1241 -3224 -1235 3152
rect -1281 -3236 -1235 -3224
rect -23 3152 23 3164
rect -23 -3224 -17 3152
rect 17 -3224 23 3152
rect -23 -3236 23 -3224
rect 1235 3152 1281 3164
rect 1235 -3224 1241 3152
rect 1275 -3224 1281 3152
rect 1235 -3236 1281 -3224
rect 2493 3152 2539 3164
rect 2493 -3224 2499 3152
rect 2533 -3224 2539 3152
rect 2493 -3236 2539 -3224
rect 3751 3152 3797 3164
rect 3751 -3224 3757 3152
rect 3791 -3224 3797 3152
rect 3751 -3236 3797 -3224
<< properties >>
string FIXED_BBOX -3908 -3367 3908 3367
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 6.0 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
