magic
tech sky130B
magscale 1 2
timestamp 1667223724
<< nwell >>
rect -3374 -3462 3374 3462
<< mvpmos >>
rect -3116 -3236 -1916 3164
rect -1858 -3236 -658 3164
rect -600 -3236 600 3164
rect 658 -3236 1858 3164
rect 1916 -3236 3116 3164
<< mvpdiff >>
rect -3174 3152 -3116 3164
rect -3174 -3224 -3162 3152
rect -3128 -3224 -3116 3152
rect -3174 -3236 -3116 -3224
rect -1916 3152 -1858 3164
rect -1916 -3224 -1904 3152
rect -1870 -3224 -1858 3152
rect -1916 -3236 -1858 -3224
rect -658 3152 -600 3164
rect -658 -3224 -646 3152
rect -612 -3224 -600 3152
rect -658 -3236 -600 -3224
rect 600 3152 658 3164
rect 600 -3224 612 3152
rect 646 -3224 658 3152
rect 600 -3236 658 -3224
rect 1858 3152 1916 3164
rect 1858 -3224 1870 3152
rect 1904 -3224 1916 3152
rect 1858 -3236 1916 -3224
rect 3116 3152 3174 3164
rect 3116 -3224 3128 3152
rect 3162 -3224 3174 3152
rect 3116 -3236 3174 -3224
<< mvpdiffc >>
rect -3162 -3224 -3128 3152
rect -1904 -3224 -1870 3152
rect -646 -3224 -612 3152
rect 612 -3224 646 3152
rect 1870 -3224 1904 3152
rect 3128 -3224 3162 3152
<< mvnsubdiff >>
rect -3308 3384 3308 3396
rect -3308 3350 -3200 3384
rect 3200 3350 3308 3384
rect -3308 3338 3308 3350
rect -3308 3288 -3250 3338
rect -3308 -3288 -3296 3288
rect -3262 -3288 -3250 3288
rect 3250 3288 3308 3338
rect -3308 -3338 -3250 -3288
rect 3250 -3288 3262 3288
rect 3296 -3288 3308 3288
rect 3250 -3338 3308 -3288
rect -3308 -3350 3308 -3338
rect -3308 -3384 -3200 -3350
rect 3200 -3384 3308 -3350
rect -3308 -3396 3308 -3384
<< mvnsubdiffcont >>
rect -3200 3350 3200 3384
rect -3296 -3288 -3262 3288
rect 3262 -3288 3296 3288
rect -3200 -3384 3200 -3350
<< poly >>
rect -3116 3245 -1916 3261
rect -3116 3211 -3100 3245
rect -1932 3211 -1916 3245
rect -3116 3164 -1916 3211
rect -1858 3245 -658 3261
rect -1858 3211 -1842 3245
rect -674 3211 -658 3245
rect -1858 3164 -658 3211
rect -600 3245 600 3261
rect -600 3211 -584 3245
rect 584 3211 600 3245
rect -600 3164 600 3211
rect 658 3245 1858 3261
rect 658 3211 674 3245
rect 1842 3211 1858 3245
rect 658 3164 1858 3211
rect 1916 3245 3116 3261
rect 1916 3211 1932 3245
rect 3100 3211 3116 3245
rect 1916 3164 3116 3211
rect -3116 -3262 -1916 -3236
rect -1858 -3262 -658 -3236
rect -600 -3262 600 -3236
rect 658 -3262 1858 -3236
rect 1916 -3262 3116 -3236
<< polycont >>
rect -3100 3211 -1932 3245
rect -1842 3211 -674 3245
rect -584 3211 584 3245
rect 674 3211 1842 3245
rect 1932 3211 3100 3245
<< locali >>
rect -3296 3350 -3200 3384
rect 3200 3350 3296 3384
rect -3296 3288 -3262 3350
rect 3262 3288 3296 3350
rect -3116 3211 -3100 3245
rect -1932 3211 -1916 3245
rect -1858 3211 -1842 3245
rect -674 3211 -658 3245
rect -600 3211 -584 3245
rect 584 3211 600 3245
rect 658 3211 674 3245
rect 1842 3211 1858 3245
rect 1916 3211 1932 3245
rect 3100 3211 3116 3245
rect -3162 3152 -3128 3168
rect -3162 -3240 -3128 -3224
rect -1904 3152 -1870 3168
rect -1904 -3240 -1870 -3224
rect -646 3152 -612 3168
rect -646 -3240 -612 -3224
rect 612 3152 646 3168
rect 612 -3240 646 -3224
rect 1870 3152 1904 3168
rect 1870 -3240 1904 -3224
rect 3128 3152 3162 3168
rect 3128 -3240 3162 -3224
rect -3296 -3350 -3262 -3288
rect 3262 -3350 3296 -3288
rect -3296 -3384 -3200 -3350
rect 3200 -3384 3296 -3350
<< viali >>
rect -3100 3211 -1932 3245
rect -1842 3211 -674 3245
rect -584 3211 584 3245
rect 674 3211 1842 3245
rect 1932 3211 3100 3245
rect -3162 -3224 -3128 3152
rect -1904 -3224 -1870 3152
rect -646 -3224 -612 3152
rect 612 -3224 646 3152
rect 1870 -3224 1904 3152
rect 3128 -3224 3162 3152
<< metal1 >>
rect -3112 3245 -1920 3251
rect -3112 3211 -3100 3245
rect -1932 3211 -1920 3245
rect -3112 3205 -1920 3211
rect -1854 3245 -662 3251
rect -1854 3211 -1842 3245
rect -674 3211 -662 3245
rect -1854 3205 -662 3211
rect -596 3245 596 3251
rect -596 3211 -584 3245
rect 584 3211 596 3245
rect -596 3205 596 3211
rect 662 3245 1854 3251
rect 662 3211 674 3245
rect 1842 3211 1854 3245
rect 662 3205 1854 3211
rect 1920 3245 3112 3251
rect 1920 3211 1932 3245
rect 3100 3211 3112 3245
rect 1920 3205 3112 3211
rect -3168 3152 -3122 3164
rect -3168 -3224 -3162 3152
rect -3128 -3224 -3122 3152
rect -3168 -3236 -3122 -3224
rect -1910 3152 -1864 3164
rect -1910 -3224 -1904 3152
rect -1870 -3224 -1864 3152
rect -1910 -3236 -1864 -3224
rect -652 3152 -606 3164
rect -652 -3224 -646 3152
rect -612 -3224 -606 3152
rect -652 -3236 -606 -3224
rect 606 3152 652 3164
rect 606 -3224 612 3152
rect 646 -3224 652 3152
rect 606 -3236 652 -3224
rect 1864 3152 1910 3164
rect 1864 -3224 1870 3152
rect 1904 -3224 1910 3152
rect 1864 -3236 1910 -3224
rect 3122 3152 3168 3164
rect 3122 -3224 3128 3152
rect 3162 -3224 3168 3152
rect 3122 -3236 3168 -3224
<< properties >>
string FIXED_BBOX -3279 -3367 3279 3367
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 6.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
