magic
tech sky130B
magscale 1 2
timestamp 1667069824
<< pwell >>
rect -3344 -5027 3344 5027
<< mvnmos >>
rect -3116 -4831 -1916 4769
rect -1858 -4831 -658 4769
rect -600 -4831 600 4769
rect 658 -4831 1858 4769
rect 1916 -4831 3116 4769
<< mvndiff >>
rect -3174 4757 -3116 4769
rect -3174 -4819 -3162 4757
rect -3128 -4819 -3116 4757
rect -3174 -4831 -3116 -4819
rect -1916 4757 -1858 4769
rect -1916 -4819 -1904 4757
rect -1870 -4819 -1858 4757
rect -1916 -4831 -1858 -4819
rect -658 4757 -600 4769
rect -658 -4819 -646 4757
rect -612 -4819 -600 4757
rect -658 -4831 -600 -4819
rect 600 4757 658 4769
rect 600 -4819 612 4757
rect 646 -4819 658 4757
rect 600 -4831 658 -4819
rect 1858 4757 1916 4769
rect 1858 -4819 1870 4757
rect 1904 -4819 1916 4757
rect 1858 -4831 1916 -4819
rect 3116 4757 3174 4769
rect 3116 -4819 3128 4757
rect 3162 -4819 3174 4757
rect 3116 -4831 3174 -4819
<< mvndiffc >>
rect -3162 -4819 -3128 4757
rect -1904 -4819 -1870 4757
rect -646 -4819 -612 4757
rect 612 -4819 646 4757
rect 1870 -4819 1904 4757
rect 3128 -4819 3162 4757
<< mvpsubdiff >>
rect -3308 4979 3308 4991
rect -3308 4945 -3200 4979
rect 3200 4945 3308 4979
rect -3308 4933 3308 4945
rect -3308 4883 -3250 4933
rect -3308 -4883 -3296 4883
rect -3262 -4883 -3250 4883
rect 3250 4883 3308 4933
rect -3308 -4933 -3250 -4883
rect 3250 -4883 3262 4883
rect 3296 -4883 3308 4883
rect 3250 -4933 3308 -4883
rect -3308 -4945 3308 -4933
rect -3308 -4979 -3200 -4945
rect 3200 -4979 3308 -4945
rect -3308 -4991 3308 -4979
<< mvpsubdiffcont >>
rect -3200 4945 3200 4979
rect -3296 -4883 -3262 4883
rect 3262 -4883 3296 4883
rect -3200 -4979 3200 -4945
<< poly >>
rect -3116 4841 -1916 4857
rect -3116 4807 -3100 4841
rect -1932 4807 -1916 4841
rect -3116 4769 -1916 4807
rect -1858 4841 -658 4857
rect -1858 4807 -1842 4841
rect -674 4807 -658 4841
rect -1858 4769 -658 4807
rect -600 4841 600 4857
rect -600 4807 -584 4841
rect 584 4807 600 4841
rect -600 4769 600 4807
rect 658 4841 1858 4857
rect 658 4807 674 4841
rect 1842 4807 1858 4841
rect 658 4769 1858 4807
rect 1916 4841 3116 4857
rect 1916 4807 1932 4841
rect 3100 4807 3116 4841
rect 1916 4769 3116 4807
rect -3116 -4857 -1916 -4831
rect -1858 -4857 -658 -4831
rect -600 -4857 600 -4831
rect 658 -4857 1858 -4831
rect 1916 -4857 3116 -4831
<< polycont >>
rect -3100 4807 -1932 4841
rect -1842 4807 -674 4841
rect -584 4807 584 4841
rect 674 4807 1842 4841
rect 1932 4807 3100 4841
<< locali >>
rect -3296 4945 -3200 4979
rect 3200 4945 3296 4979
rect -3296 4883 -3262 4945
rect 3262 4883 3296 4945
rect -3116 4807 -3100 4841
rect -1932 4807 -1916 4841
rect -1858 4807 -1842 4841
rect -674 4807 -658 4841
rect -600 4807 -584 4841
rect 584 4807 600 4841
rect 658 4807 674 4841
rect 1842 4807 1858 4841
rect 1916 4807 1932 4841
rect 3100 4807 3116 4841
rect -3162 4757 -3128 4773
rect -3162 -4835 -3128 -4819
rect -1904 4757 -1870 4773
rect -1904 -4835 -1870 -4819
rect -646 4757 -612 4773
rect -646 -4835 -612 -4819
rect 612 4757 646 4773
rect 612 -4835 646 -4819
rect 1870 4757 1904 4773
rect 1870 -4835 1904 -4819
rect 3128 4757 3162 4773
rect 3128 -4835 3162 -4819
rect -3296 -4945 -3262 -4883
rect 3262 -4945 3296 -4883
rect -3296 -4979 -3200 -4945
rect 3200 -4979 3296 -4945
<< viali >>
rect -3100 4807 -1932 4841
rect -1842 4807 -674 4841
rect -584 4807 584 4841
rect 674 4807 1842 4841
rect 1932 4807 3100 4841
rect -3162 -4819 -3128 4757
rect -1904 -4819 -1870 4757
rect -646 -4819 -612 4757
rect 612 -4819 646 4757
rect 1870 -4819 1904 4757
rect 3128 -4819 3162 4757
<< metal1 >>
rect -3112 4841 -1920 4847
rect -3112 4807 -3100 4841
rect -1932 4807 -1920 4841
rect -3112 4801 -1920 4807
rect -1854 4841 -662 4847
rect -1854 4807 -1842 4841
rect -674 4807 -662 4841
rect -1854 4801 -662 4807
rect -596 4841 596 4847
rect -596 4807 -584 4841
rect 584 4807 596 4841
rect -596 4801 596 4807
rect 662 4841 1854 4847
rect 662 4807 674 4841
rect 1842 4807 1854 4841
rect 662 4801 1854 4807
rect 1920 4841 3112 4847
rect 1920 4807 1932 4841
rect 3100 4807 3112 4841
rect 1920 4801 3112 4807
rect -3168 4757 -3122 4769
rect -3168 -4819 -3162 4757
rect -3128 -4819 -3122 4757
rect -3168 -4831 -3122 -4819
rect -1910 4757 -1864 4769
rect -1910 -4819 -1904 4757
rect -1870 -4819 -1864 4757
rect -1910 -4831 -1864 -4819
rect -652 4757 -606 4769
rect -652 -4819 -646 4757
rect -612 -4819 -606 4757
rect -652 -4831 -606 -4819
rect 606 4757 652 4769
rect 606 -4819 612 4757
rect 646 -4819 652 4757
rect 606 -4831 652 -4819
rect 1864 4757 1910 4769
rect 1864 -4819 1870 4757
rect 1904 -4819 1910 4757
rect 1864 -4831 1910 -4819
rect 3122 4757 3168 4769
rect 3122 -4819 3128 4757
rect 3162 -4819 3168 4757
rect 3122 -4831 3168 -4819
<< properties >>
string FIXED_BBOX -3279 -4962 3279 4962
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 48.0 l 6.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
