magic
tech sky130B
magscale 1 2
timestamp 1667934541
<< pwell >>
rect -3344 -5027 3344 5027
<< mvnmos >>
rect -3116 -4831 -1916 4769
rect -1858 -4831 -658 4769
rect -600 -4831 600 4769
rect 658 -4831 1858 4769
rect 1916 -4831 3116 4769
<< mvndiff >>
rect -3174 3799 -3116 4769
rect -3174 -3861 -3162 3799
rect -3128 -3861 -3116 3799
rect -3174 -4831 -3116 -3861
rect -1916 3799 -1858 4769
rect -1916 -3861 -1904 3799
rect -1870 -3861 -1858 3799
rect -1916 -4831 -1858 -3861
rect -658 3799 -600 4769
rect -658 -3861 -646 3799
rect -612 -3861 -600 3799
rect -658 -4831 -600 -3861
rect 600 3799 658 4769
rect 600 -3861 612 3799
rect 646 -3861 658 3799
rect 600 -4831 658 -3861
rect 1858 3799 1916 4769
rect 1858 -3861 1870 3799
rect 1904 -3861 1916 3799
rect 1858 -4831 1916 -3861
rect 3116 3799 3174 4769
rect 3116 -3861 3128 3799
rect 3162 -3861 3174 3799
rect 3116 -4831 3174 -3861
<< mvndiffc >>
rect -3162 -3861 -3128 3799
rect -1904 -3861 -1870 3799
rect -646 -3861 -612 3799
rect 612 -3861 646 3799
rect 1870 -3861 1904 3799
rect 3128 -3861 3162 3799
<< mvpsubdiff >>
rect -3308 4933 3308 4991
rect -3308 -4933 -3250 4933
rect 3250 -4933 3308 4933
rect -3308 -4945 3308 -4933
rect -3308 -4979 -2560 -4945
rect 2560 -4979 3308 -4945
rect -3308 -4991 3308 -4979
<< mvpsubdiffcont >>
rect -2560 -4979 2560 -4945
<< poly >>
rect -3058 4841 -1974 4857
rect -3058 4824 -3042 4841
rect -3116 4807 -3042 4824
rect -1990 4824 -1974 4841
rect -1800 4841 -716 4857
rect -1800 4824 -1784 4841
rect -1990 4807 -1916 4824
rect -3116 4769 -1916 4807
rect -1858 4807 -1784 4824
rect -732 4824 -716 4841
rect -542 4841 542 4857
rect -542 4824 -526 4841
rect -732 4807 -658 4824
rect -1858 4769 -658 4807
rect -600 4807 -526 4824
rect 526 4824 542 4841
rect 716 4841 1800 4857
rect 716 4824 732 4841
rect 526 4807 600 4824
rect -600 4769 600 4807
rect 658 4807 732 4824
rect 1784 4824 1800 4841
rect 1974 4841 3058 4857
rect 1974 4824 1990 4841
rect 1784 4807 1858 4824
rect 658 4769 1858 4807
rect 1916 4807 1990 4824
rect 3042 4824 3058 4841
rect 3042 4807 3116 4824
rect 1916 4769 3116 4807
rect -3116 -4857 -1916 -4831
rect -1858 -4857 -658 -4831
rect -600 -4857 600 -4831
rect 658 -4857 1858 -4831
rect 1916 -4857 3116 -4831
<< polycont >>
rect -3042 4807 -1990 4841
rect -1784 4807 -732 4841
rect -526 4807 526 4841
rect 732 4807 1784 4841
rect 1990 4807 3042 4841
<< locali >>
rect -3058 4807 -3042 4841
rect -1990 4807 -1974 4841
rect -1800 4807 -1784 4841
rect -732 4807 -716 4841
rect -542 4807 -526 4841
rect 526 4807 542 4841
rect 716 4807 732 4841
rect 1784 4807 1800 4841
rect 1974 4807 1990 4841
rect 3042 4807 3058 4841
rect -3162 3799 -3128 3815
rect -3162 -3877 -3128 -3861
rect -1904 3799 -1870 3815
rect -1904 -3877 -1870 -3861
rect -646 3799 -612 3815
rect -646 -3877 -612 -3861
rect 612 3799 646 3815
rect 612 -3877 646 -3861
rect 1870 3799 1904 3815
rect 1870 -3877 1904 -3861
rect 3128 3799 3162 3815
rect 3128 -3877 3162 -3861
rect -2576 -4979 -2560 -4945
rect 2560 -4979 2576 -4945
<< viali >>
rect -3042 4807 -1990 4841
rect -1784 4807 -732 4841
rect -526 4807 526 4841
rect 732 4807 1784 4841
rect 1990 4807 3042 4841
rect -3162 -3861 -3128 3799
rect -1904 -3861 -1870 3799
rect -646 -3861 -612 3799
rect 612 -3861 646 3799
rect 1870 -3861 1904 3799
rect 3128 -3861 3162 3799
<< metal1 >>
rect -3054 4841 -1978 4847
rect -3054 4807 -3042 4841
rect -1990 4807 -1978 4841
rect -3054 4801 -1978 4807
rect -1796 4841 -720 4847
rect -1796 4807 -1784 4841
rect -732 4807 -720 4841
rect -1796 4801 -720 4807
rect -538 4841 538 4847
rect -538 4807 -526 4841
rect 526 4807 538 4841
rect -538 4801 538 4807
rect 720 4841 1796 4847
rect 720 4807 732 4841
rect 1784 4807 1796 4841
rect 720 4801 1796 4807
rect 1978 4841 3054 4847
rect 1978 4807 1990 4841
rect 3042 4807 3054 4841
rect 1978 4801 3054 4807
rect -3168 3799 -3122 3811
rect -3168 -3861 -3162 3799
rect -3128 -3861 -3122 3799
rect -3168 -3873 -3122 -3861
rect -1910 3799 -1864 3811
rect -1910 -3861 -1904 3799
rect -1870 -3861 -1864 3799
rect -1910 -3873 -1864 -3861
rect -652 3799 -606 3811
rect -652 -3861 -646 3799
rect -612 -3861 -606 3799
rect -652 -3873 -606 -3861
rect 606 3799 652 3811
rect 606 -3861 612 3799
rect 646 -3861 652 3799
rect 606 -3873 652 -3861
rect 1864 3799 1910 3811
rect 1864 -3861 1870 3799
rect 1904 -3861 1910 3799
rect 1864 -3873 1910 -3861
rect 3122 3799 3168 3811
rect 3122 -3861 3128 3799
rect 3162 -3861 3168 3799
rect 3122 -3873 3168 -3861
<< properties >>
string FIXED_BBOX -3279 -4962 3279 4962
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 48.0 l 6.0 m 1 nf 5 diffcov 80 polycov 90 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 80 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 80 viadrn 80 viagate 90 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
