magic
tech sky130B
magscale 1 2
timestamp 1667069824
<< nwell >>
rect -2745 -10109 2745 10109
<< mvpmos >>
rect -2487 5012 -1287 9812
rect -1229 5012 -29 9812
rect 29 5012 1229 9812
rect 1287 5012 2487 9812
rect -2487 47 -1287 4847
rect -1229 47 -29 4847
rect 29 47 1229 4847
rect 1287 47 2487 4847
rect -2487 -4918 -1287 -118
rect -1229 -4918 -29 -118
rect 29 -4918 1229 -118
rect 1287 -4918 2487 -118
rect -2487 -9883 -1287 -5083
rect -1229 -9883 -29 -5083
rect 29 -9883 1229 -5083
rect 1287 -9883 2487 -5083
<< mvpdiff >>
rect -2545 9800 -2487 9812
rect -2545 5024 -2533 9800
rect -2499 5024 -2487 9800
rect -2545 5012 -2487 5024
rect -1287 9800 -1229 9812
rect -1287 5024 -1275 9800
rect -1241 5024 -1229 9800
rect -1287 5012 -1229 5024
rect -29 9800 29 9812
rect -29 5024 -17 9800
rect 17 5024 29 9800
rect -29 5012 29 5024
rect 1229 9800 1287 9812
rect 1229 5024 1241 9800
rect 1275 5024 1287 9800
rect 1229 5012 1287 5024
rect 2487 9800 2545 9812
rect 2487 5024 2499 9800
rect 2533 5024 2545 9800
rect 2487 5012 2545 5024
rect -2545 4835 -2487 4847
rect -2545 59 -2533 4835
rect -2499 59 -2487 4835
rect -2545 47 -2487 59
rect -1287 4835 -1229 4847
rect -1287 59 -1275 4835
rect -1241 59 -1229 4835
rect -1287 47 -1229 59
rect -29 4835 29 4847
rect -29 59 -17 4835
rect 17 59 29 4835
rect -29 47 29 59
rect 1229 4835 1287 4847
rect 1229 59 1241 4835
rect 1275 59 1287 4835
rect 1229 47 1287 59
rect 2487 4835 2545 4847
rect 2487 59 2499 4835
rect 2533 59 2545 4835
rect 2487 47 2545 59
rect -2545 -130 -2487 -118
rect -2545 -4906 -2533 -130
rect -2499 -4906 -2487 -130
rect -2545 -4918 -2487 -4906
rect -1287 -130 -1229 -118
rect -1287 -4906 -1275 -130
rect -1241 -4906 -1229 -130
rect -1287 -4918 -1229 -4906
rect -29 -130 29 -118
rect -29 -4906 -17 -130
rect 17 -4906 29 -130
rect -29 -4918 29 -4906
rect 1229 -130 1287 -118
rect 1229 -4906 1241 -130
rect 1275 -4906 1287 -130
rect 1229 -4918 1287 -4906
rect 2487 -130 2545 -118
rect 2487 -4906 2499 -130
rect 2533 -4906 2545 -130
rect 2487 -4918 2545 -4906
rect -2545 -5095 -2487 -5083
rect -2545 -9871 -2533 -5095
rect -2499 -9871 -2487 -5095
rect -2545 -9883 -2487 -9871
rect -1287 -5095 -1229 -5083
rect -1287 -9871 -1275 -5095
rect -1241 -9871 -1229 -5095
rect -1287 -9883 -1229 -9871
rect -29 -5095 29 -5083
rect -29 -9871 -17 -5095
rect 17 -9871 29 -5095
rect -29 -9883 29 -9871
rect 1229 -5095 1287 -5083
rect 1229 -9871 1241 -5095
rect 1275 -9871 1287 -5095
rect 1229 -9883 1287 -9871
rect 2487 -5095 2545 -5083
rect 2487 -9871 2499 -5095
rect 2533 -9871 2545 -5095
rect 2487 -9883 2545 -9871
<< mvpdiffc >>
rect -2533 5024 -2499 9800
rect -1275 5024 -1241 9800
rect -17 5024 17 9800
rect 1241 5024 1275 9800
rect 2499 5024 2533 9800
rect -2533 59 -2499 4835
rect -1275 59 -1241 4835
rect -17 59 17 4835
rect 1241 59 1275 4835
rect 2499 59 2533 4835
rect -2533 -4906 -2499 -130
rect -1275 -4906 -1241 -130
rect -17 -4906 17 -130
rect 1241 -4906 1275 -130
rect 2499 -4906 2533 -130
rect -2533 -9871 -2499 -5095
rect -1275 -9871 -1241 -5095
rect -17 -9871 17 -5095
rect 1241 -9871 1275 -5095
rect 2499 -9871 2533 -5095
<< mvnsubdiff >>
rect -2679 10031 2679 10043
rect -2679 9997 -2571 10031
rect 2571 9997 2679 10031
rect -2679 9985 2679 9997
rect -2679 9935 -2621 9985
rect -2679 -9935 -2667 9935
rect -2633 -9935 -2621 9935
rect 2621 9935 2679 9985
rect -2679 -9985 -2621 -9935
rect 2621 -9935 2633 9935
rect 2667 -9935 2679 9935
rect 2621 -9985 2679 -9935
rect -2679 -9997 2679 -9985
rect -2679 -10031 -2571 -9997
rect 2571 -10031 2679 -9997
rect -2679 -10043 2679 -10031
<< mvnsubdiffcont >>
rect -2571 9997 2571 10031
rect -2667 -9935 -2633 9935
rect 2633 -9935 2667 9935
rect -2571 -10031 2571 -9997
<< poly >>
rect -2487 9893 -1287 9909
rect -2487 9859 -2471 9893
rect -1303 9859 -1287 9893
rect -2487 9812 -1287 9859
rect -1229 9893 -29 9909
rect -1229 9859 -1213 9893
rect -45 9859 -29 9893
rect -1229 9812 -29 9859
rect 29 9893 1229 9909
rect 29 9859 45 9893
rect 1213 9859 1229 9893
rect 29 9812 1229 9859
rect 1287 9893 2487 9909
rect 1287 9859 1303 9893
rect 2471 9859 2487 9893
rect 1287 9812 2487 9859
rect -2487 4986 -1287 5012
rect -1229 4986 -29 5012
rect 29 4986 1229 5012
rect 1287 4986 2487 5012
rect -2487 4928 -1287 4944
rect -2487 4894 -2471 4928
rect -1303 4894 -1287 4928
rect -2487 4847 -1287 4894
rect -1229 4928 -29 4944
rect -1229 4894 -1213 4928
rect -45 4894 -29 4928
rect -1229 4847 -29 4894
rect 29 4928 1229 4944
rect 29 4894 45 4928
rect 1213 4894 1229 4928
rect 29 4847 1229 4894
rect 1287 4928 2487 4944
rect 1287 4894 1303 4928
rect 2471 4894 2487 4928
rect 1287 4847 2487 4894
rect -2487 21 -1287 47
rect -1229 21 -29 47
rect 29 21 1229 47
rect 1287 21 2487 47
rect -2487 -37 -1287 -21
rect -2487 -71 -2471 -37
rect -1303 -71 -1287 -37
rect -2487 -118 -1287 -71
rect -1229 -37 -29 -21
rect -1229 -71 -1213 -37
rect -45 -71 -29 -37
rect -1229 -118 -29 -71
rect 29 -37 1229 -21
rect 29 -71 45 -37
rect 1213 -71 1229 -37
rect 29 -118 1229 -71
rect 1287 -37 2487 -21
rect 1287 -71 1303 -37
rect 2471 -71 2487 -37
rect 1287 -118 2487 -71
rect -2487 -4944 -1287 -4918
rect -1229 -4944 -29 -4918
rect 29 -4944 1229 -4918
rect 1287 -4944 2487 -4918
rect -2487 -5002 -1287 -4986
rect -2487 -5036 -2471 -5002
rect -1303 -5036 -1287 -5002
rect -2487 -5083 -1287 -5036
rect -1229 -5002 -29 -4986
rect -1229 -5036 -1213 -5002
rect -45 -5036 -29 -5002
rect -1229 -5083 -29 -5036
rect 29 -5002 1229 -4986
rect 29 -5036 45 -5002
rect 1213 -5036 1229 -5002
rect 29 -5083 1229 -5036
rect 1287 -5002 2487 -4986
rect 1287 -5036 1303 -5002
rect 2471 -5036 2487 -5002
rect 1287 -5083 2487 -5036
rect -2487 -9909 -1287 -9883
rect -1229 -9909 -29 -9883
rect 29 -9909 1229 -9883
rect 1287 -9909 2487 -9883
<< polycont >>
rect -2471 9859 -1303 9893
rect -1213 9859 -45 9893
rect 45 9859 1213 9893
rect 1303 9859 2471 9893
rect -2471 4894 -1303 4928
rect -1213 4894 -45 4928
rect 45 4894 1213 4928
rect 1303 4894 2471 4928
rect -2471 -71 -1303 -37
rect -1213 -71 -45 -37
rect 45 -71 1213 -37
rect 1303 -71 2471 -37
rect -2471 -5036 -1303 -5002
rect -1213 -5036 -45 -5002
rect 45 -5036 1213 -5002
rect 1303 -5036 2471 -5002
<< locali >>
rect -2667 9997 -2571 10031
rect 2571 9997 2667 10031
rect -2667 9935 -2633 9997
rect 2633 9935 2667 9997
rect -2487 9859 -2471 9893
rect -1303 9859 -1287 9893
rect -1229 9859 -1213 9893
rect -45 9859 -29 9893
rect 29 9859 45 9893
rect 1213 9859 1229 9893
rect 1287 9859 1303 9893
rect 2471 9859 2487 9893
rect -2533 9800 -2499 9816
rect -2533 5008 -2499 5024
rect -1275 9800 -1241 9816
rect -1275 5008 -1241 5024
rect -17 9800 17 9816
rect -17 5008 17 5024
rect 1241 9800 1275 9816
rect 1241 5008 1275 5024
rect 2499 9800 2533 9816
rect 2499 5008 2533 5024
rect -2487 4894 -2471 4928
rect -1303 4894 -1287 4928
rect -1229 4894 -1213 4928
rect -45 4894 -29 4928
rect 29 4894 45 4928
rect 1213 4894 1229 4928
rect 1287 4894 1303 4928
rect 2471 4894 2487 4928
rect -2533 4835 -2499 4851
rect -2533 43 -2499 59
rect -1275 4835 -1241 4851
rect -1275 43 -1241 59
rect -17 4835 17 4851
rect -17 43 17 59
rect 1241 4835 1275 4851
rect 1241 43 1275 59
rect 2499 4835 2533 4851
rect 2499 43 2533 59
rect -2487 -71 -2471 -37
rect -1303 -71 -1287 -37
rect -1229 -71 -1213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1213 -71 1229 -37
rect 1287 -71 1303 -37
rect 2471 -71 2487 -37
rect -2533 -130 -2499 -114
rect -2533 -4922 -2499 -4906
rect -1275 -130 -1241 -114
rect -1275 -4922 -1241 -4906
rect -17 -130 17 -114
rect -17 -4922 17 -4906
rect 1241 -130 1275 -114
rect 1241 -4922 1275 -4906
rect 2499 -130 2533 -114
rect 2499 -4922 2533 -4906
rect -2487 -5036 -2471 -5002
rect -1303 -5036 -1287 -5002
rect -1229 -5036 -1213 -5002
rect -45 -5036 -29 -5002
rect 29 -5036 45 -5002
rect 1213 -5036 1229 -5002
rect 1287 -5036 1303 -5002
rect 2471 -5036 2487 -5002
rect -2533 -5095 -2499 -5079
rect -2533 -9887 -2499 -9871
rect -1275 -5095 -1241 -5079
rect -1275 -9887 -1241 -9871
rect -17 -5095 17 -5079
rect -17 -9887 17 -9871
rect 1241 -5095 1275 -5079
rect 1241 -9887 1275 -9871
rect 2499 -5095 2533 -5079
rect 2499 -9887 2533 -9871
rect -2667 -9997 -2633 -9935
rect 2633 -9997 2667 -9935
rect -2667 -10031 -2571 -9997
rect 2571 -10031 2667 -9997
<< viali >>
rect -2471 9859 -1303 9893
rect -1213 9859 -45 9893
rect 45 9859 1213 9893
rect 1303 9859 2471 9893
rect -2533 5024 -2499 9800
rect -1275 5024 -1241 9800
rect -17 5024 17 9800
rect 1241 5024 1275 9800
rect 2499 5024 2533 9800
rect -2471 4894 -1303 4928
rect -1213 4894 -45 4928
rect 45 4894 1213 4928
rect 1303 4894 2471 4928
rect -2533 59 -2499 4835
rect -1275 59 -1241 4835
rect -17 59 17 4835
rect 1241 59 1275 4835
rect 2499 59 2533 4835
rect -2471 -71 -1303 -37
rect -1213 -71 -45 -37
rect 45 -71 1213 -37
rect 1303 -71 2471 -37
rect -2533 -4906 -2499 -130
rect -1275 -4906 -1241 -130
rect -17 -4906 17 -130
rect 1241 -4906 1275 -130
rect 2499 -4906 2533 -130
rect -2471 -5036 -1303 -5002
rect -1213 -5036 -45 -5002
rect 45 -5036 1213 -5002
rect 1303 -5036 2471 -5002
rect -2533 -9871 -2499 -5095
rect -1275 -9871 -1241 -5095
rect -17 -9871 17 -5095
rect 1241 -9871 1275 -5095
rect 2499 -9871 2533 -5095
<< metal1 >>
rect -2483 9893 -1291 9899
rect -2483 9859 -2471 9893
rect -1303 9859 -1291 9893
rect -2483 9853 -1291 9859
rect -1225 9893 -33 9899
rect -1225 9859 -1213 9893
rect -45 9859 -33 9893
rect -1225 9853 -33 9859
rect 33 9893 1225 9899
rect 33 9859 45 9893
rect 1213 9859 1225 9893
rect 33 9853 1225 9859
rect 1291 9893 2483 9899
rect 1291 9859 1303 9893
rect 2471 9859 2483 9893
rect 1291 9853 2483 9859
rect -2539 9800 -2493 9812
rect -2539 5024 -2533 9800
rect -2499 5024 -2493 9800
rect -2539 5012 -2493 5024
rect -1281 9800 -1235 9812
rect -1281 5024 -1275 9800
rect -1241 5024 -1235 9800
rect -1281 5012 -1235 5024
rect -23 9800 23 9812
rect -23 5024 -17 9800
rect 17 5024 23 9800
rect -23 5012 23 5024
rect 1235 9800 1281 9812
rect 1235 5024 1241 9800
rect 1275 5024 1281 9800
rect 1235 5012 1281 5024
rect 2493 9800 2539 9812
rect 2493 5024 2499 9800
rect 2533 5024 2539 9800
rect 2493 5012 2539 5024
rect -2483 4928 -1291 4934
rect -2483 4894 -2471 4928
rect -1303 4894 -1291 4928
rect -2483 4888 -1291 4894
rect -1225 4928 -33 4934
rect -1225 4894 -1213 4928
rect -45 4894 -33 4928
rect -1225 4888 -33 4894
rect 33 4928 1225 4934
rect 33 4894 45 4928
rect 1213 4894 1225 4928
rect 33 4888 1225 4894
rect 1291 4928 2483 4934
rect 1291 4894 1303 4928
rect 2471 4894 2483 4928
rect 1291 4888 2483 4894
rect -2539 4835 -2493 4847
rect -2539 59 -2533 4835
rect -2499 59 -2493 4835
rect -2539 47 -2493 59
rect -1281 4835 -1235 4847
rect -1281 59 -1275 4835
rect -1241 59 -1235 4835
rect -1281 47 -1235 59
rect -23 4835 23 4847
rect -23 59 -17 4835
rect 17 59 23 4835
rect -23 47 23 59
rect 1235 4835 1281 4847
rect 1235 59 1241 4835
rect 1275 59 1281 4835
rect 1235 47 1281 59
rect 2493 4835 2539 4847
rect 2493 59 2499 4835
rect 2533 59 2539 4835
rect 2493 47 2539 59
rect -2483 -37 -1291 -31
rect -2483 -71 -2471 -37
rect -1303 -71 -1291 -37
rect -2483 -77 -1291 -71
rect -1225 -37 -33 -31
rect -1225 -71 -1213 -37
rect -45 -71 -33 -37
rect -1225 -77 -33 -71
rect 33 -37 1225 -31
rect 33 -71 45 -37
rect 1213 -71 1225 -37
rect 33 -77 1225 -71
rect 1291 -37 2483 -31
rect 1291 -71 1303 -37
rect 2471 -71 2483 -37
rect 1291 -77 2483 -71
rect -2539 -130 -2493 -118
rect -2539 -4906 -2533 -130
rect -2499 -4906 -2493 -130
rect -2539 -4918 -2493 -4906
rect -1281 -130 -1235 -118
rect -1281 -4906 -1275 -130
rect -1241 -4906 -1235 -130
rect -1281 -4918 -1235 -4906
rect -23 -130 23 -118
rect -23 -4906 -17 -130
rect 17 -4906 23 -130
rect -23 -4918 23 -4906
rect 1235 -130 1281 -118
rect 1235 -4906 1241 -130
rect 1275 -4906 1281 -130
rect 1235 -4918 1281 -4906
rect 2493 -130 2539 -118
rect 2493 -4906 2499 -130
rect 2533 -4906 2539 -130
rect 2493 -4918 2539 -4906
rect -2483 -5002 -1291 -4996
rect -2483 -5036 -2471 -5002
rect -1303 -5036 -1291 -5002
rect -2483 -5042 -1291 -5036
rect -1225 -5002 -33 -4996
rect -1225 -5036 -1213 -5002
rect -45 -5036 -33 -5002
rect -1225 -5042 -33 -5036
rect 33 -5002 1225 -4996
rect 33 -5036 45 -5002
rect 1213 -5036 1225 -5002
rect 33 -5042 1225 -5036
rect 1291 -5002 2483 -4996
rect 1291 -5036 1303 -5002
rect 2471 -5036 2483 -5002
rect 1291 -5042 2483 -5036
rect -2539 -5095 -2493 -5083
rect -2539 -9871 -2533 -5095
rect -2499 -9871 -2493 -5095
rect -2539 -9883 -2493 -9871
rect -1281 -5095 -1235 -5083
rect -1281 -9871 -1275 -5095
rect -1241 -9871 -1235 -5095
rect -1281 -9883 -1235 -9871
rect -23 -5095 23 -5083
rect -23 -9871 -17 -5095
rect 17 -9871 23 -5095
rect -23 -9883 23 -9871
rect 1235 -5095 1281 -5083
rect 1235 -9871 1241 -5095
rect 1275 -9871 1281 -5095
rect 1235 -9883 1281 -9871
rect 2493 -5095 2539 -5083
rect 2493 -9871 2499 -5095
rect 2533 -9871 2539 -5095
rect 2493 -9883 2539 -9871
<< properties >>
string FIXED_BBOX -2650 -10014 2650 10014
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 24.0 l 6.0 m 4 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
