magic
tech sky130B
magscale 1 2
timestamp 1667934541
<< nwell >>
rect -2745 -2662 2745 2662
<< mvpmos >>
rect -2487 -2436 -1287 2364
rect -1229 -2436 -29 2364
rect 29 -2436 1229 2364
rect 1287 -2436 2487 2364
<< mvpdiff >>
rect -2545 1874 -2487 2364
rect -2545 -1946 -2533 1874
rect -2499 -1946 -2487 1874
rect -2545 -2436 -2487 -1946
rect -1287 1874 -1229 2364
rect -1287 -1946 -1275 1874
rect -1241 -1946 -1229 1874
rect -1287 -2436 -1229 -1946
rect -29 1874 29 2364
rect -29 -1946 -17 1874
rect 17 -1946 29 1874
rect -29 -2436 29 -1946
rect 1229 1874 1287 2364
rect 1229 -1946 1241 1874
rect 1275 -1946 1287 1874
rect 1229 -2436 1287 -1946
rect 2487 1874 2545 2364
rect 2487 -1946 2499 1874
rect 2533 -1946 2545 1874
rect 2487 -2436 2545 -1946
<< mvpdiffc >>
rect -2533 -1946 -2499 1874
rect -1275 -1946 -1241 1874
rect -17 -1946 17 1874
rect 1241 -1946 1275 1874
rect 2499 -1946 2533 1874
<< mvnsubdiff >>
rect -2679 2584 2679 2596
rect -2679 2550 -2057 2584
rect 2057 2550 2679 2584
rect -2679 2538 2679 2550
rect -2679 -2538 -2621 2538
rect 2621 -2538 2679 2538
rect -2679 -2596 2679 -2538
<< mvnsubdiffcont >>
rect -2057 2550 2057 2584
<< poly >>
rect -2429 2445 -1345 2461
rect -2429 2428 -2413 2445
rect -2487 2411 -2413 2428
rect -1361 2428 -1345 2445
rect -1171 2445 -87 2461
rect -1171 2428 -1155 2445
rect -1361 2411 -1287 2428
rect -2487 2364 -1287 2411
rect -1229 2411 -1155 2428
rect -103 2428 -87 2445
rect 87 2445 1171 2461
rect 87 2428 103 2445
rect -103 2411 -29 2428
rect -1229 2364 -29 2411
rect 29 2411 103 2428
rect 1155 2428 1171 2445
rect 1345 2445 2429 2461
rect 1345 2428 1361 2445
rect 1155 2411 1229 2428
rect 29 2364 1229 2411
rect 1287 2411 1361 2428
rect 2413 2428 2429 2445
rect 2413 2411 2487 2428
rect 1287 2364 2487 2411
rect -2487 -2462 -1287 -2436
rect -1229 -2462 -29 -2436
rect 29 -2462 1229 -2436
rect 1287 -2462 2487 -2436
<< polycont >>
rect -2413 2411 -1361 2445
rect -1155 2411 -103 2445
rect 103 2411 1155 2445
rect 1361 2411 2413 2445
<< locali >>
rect -2073 2550 -2057 2584
rect 2057 2550 2073 2584
rect -2429 2411 -2413 2445
rect -1361 2411 -1345 2445
rect -1171 2411 -1155 2445
rect -103 2411 -87 2445
rect 87 2411 103 2445
rect 1155 2411 1171 2445
rect 1345 2411 1361 2445
rect 2413 2411 2429 2445
rect -2533 1874 -2499 1890
rect -2533 -1962 -2499 -1946
rect -1275 1874 -1241 1890
rect -1275 -1962 -1241 -1946
rect -17 1874 17 1890
rect -17 -1962 17 -1946
rect 1241 1874 1275 1890
rect 1241 -1962 1275 -1946
rect 2499 1874 2533 1890
rect 2499 -1962 2533 -1946
<< viali >>
rect -2413 2411 -1361 2445
rect -1155 2411 -103 2445
rect 103 2411 1155 2445
rect 1361 2411 2413 2445
rect -2533 -1946 -2499 1874
rect -1275 -1946 -1241 1874
rect -17 -1946 17 1874
rect 1241 -1946 1275 1874
rect 2499 -1946 2533 1874
<< metal1 >>
rect -2425 2445 -1349 2451
rect -2425 2411 -2413 2445
rect -1361 2411 -1349 2445
rect -2425 2405 -1349 2411
rect -1167 2445 -91 2451
rect -1167 2411 -1155 2445
rect -103 2411 -91 2445
rect -1167 2405 -91 2411
rect 91 2445 1167 2451
rect 91 2411 103 2445
rect 1155 2411 1167 2445
rect 91 2405 1167 2411
rect 1349 2445 2425 2451
rect 1349 2411 1361 2445
rect 2413 2411 2425 2445
rect 1349 2405 2425 2411
rect -2539 1874 -2493 1886
rect -2539 -1946 -2533 1874
rect -2499 -1946 -2493 1874
rect -2539 -1958 -2493 -1946
rect -1281 1874 -1235 1886
rect -1281 -1946 -1275 1874
rect -1241 -1946 -1235 1874
rect -1281 -1958 -1235 -1946
rect -23 1874 23 1886
rect -23 -1946 -17 1874
rect 17 -1946 23 1874
rect -23 -1958 23 -1946
rect 1235 1874 1281 1886
rect 1235 -1946 1241 1874
rect 1275 -1946 1281 1874
rect 1235 -1958 1281 -1946
rect 2493 1874 2539 1886
rect 2493 -1946 2499 1874
rect 2533 -1946 2539 1874
rect 2493 -1958 2539 -1946
<< properties >>
string FIXED_BBOX -2650 -2567 2650 2567
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 24.0 l 6.0 m 1 nf 4 diffcov 80 polycov 90 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 80 rlcov 80 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 80 viadrn 80 viagate 90 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
