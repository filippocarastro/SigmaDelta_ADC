magic
tech sky130B
magscale 1 2
timestamp 1667934541
<< nwell >>
rect -10293 -2662 10293 2662
<< mvpmos >>
rect -10035 -2364 -8835 2436
rect -8777 -2364 -7577 2436
rect -7519 -2364 -6319 2436
rect -6261 -2364 -5061 2436
rect -5003 -2364 -3803 2436
rect -3745 -2364 -2545 2436
rect -2487 -2364 -1287 2436
rect -1229 -2364 -29 2436
rect 29 -2364 1229 2436
rect 1287 -2364 2487 2436
rect 2545 -2364 3745 2436
rect 3803 -2364 5003 2436
rect 5061 -2364 6261 2436
rect 6319 -2364 7519 2436
rect 7577 -2364 8777 2436
rect 8835 -2364 10035 2436
<< mvpdiff >>
rect -10093 1946 -10035 2436
rect -10093 -1874 -10081 1946
rect -10047 -1874 -10035 1946
rect -10093 -2364 -10035 -1874
rect -8835 1946 -8777 2436
rect -8835 -1874 -8823 1946
rect -8789 -1874 -8777 1946
rect -8835 -2364 -8777 -1874
rect -7577 1946 -7519 2436
rect -7577 -1874 -7565 1946
rect -7531 -1874 -7519 1946
rect -7577 -2364 -7519 -1874
rect -6319 1946 -6261 2436
rect -6319 -1874 -6307 1946
rect -6273 -1874 -6261 1946
rect -6319 -2364 -6261 -1874
rect -5061 1946 -5003 2436
rect -5061 -1874 -5049 1946
rect -5015 -1874 -5003 1946
rect -5061 -2364 -5003 -1874
rect -3803 1946 -3745 2436
rect -3803 -1874 -3791 1946
rect -3757 -1874 -3745 1946
rect -3803 -2364 -3745 -1874
rect -2545 1946 -2487 2436
rect -2545 -1874 -2533 1946
rect -2499 -1874 -2487 1946
rect -2545 -2364 -2487 -1874
rect -1287 1946 -1229 2436
rect -1287 -1874 -1275 1946
rect -1241 -1874 -1229 1946
rect -1287 -2364 -1229 -1874
rect -29 1946 29 2436
rect -29 -1874 -17 1946
rect 17 -1874 29 1946
rect -29 -2364 29 -1874
rect 1229 1946 1287 2436
rect 1229 -1874 1241 1946
rect 1275 -1874 1287 1946
rect 1229 -2364 1287 -1874
rect 2487 1946 2545 2436
rect 2487 -1874 2499 1946
rect 2533 -1874 2545 1946
rect 2487 -2364 2545 -1874
rect 3745 1946 3803 2436
rect 3745 -1874 3757 1946
rect 3791 -1874 3803 1946
rect 3745 -2364 3803 -1874
rect 5003 1946 5061 2436
rect 5003 -1874 5015 1946
rect 5049 -1874 5061 1946
rect 5003 -2364 5061 -1874
rect 6261 1946 6319 2436
rect 6261 -1874 6273 1946
rect 6307 -1874 6319 1946
rect 6261 -2364 6319 -1874
rect 7519 1946 7577 2436
rect 7519 -1874 7531 1946
rect 7565 -1874 7577 1946
rect 7519 -2364 7577 -1874
rect 8777 1946 8835 2436
rect 8777 -1874 8789 1946
rect 8823 -1874 8835 1946
rect 8777 -2364 8835 -1874
rect 10035 1946 10093 2436
rect 10035 -1874 10047 1946
rect 10081 -1874 10093 1946
rect 10035 -2364 10093 -1874
<< mvpdiffc >>
rect -10081 -1874 -10047 1946
rect -8823 -1874 -8789 1946
rect -7565 -1874 -7531 1946
rect -6307 -1874 -6273 1946
rect -5049 -1874 -5015 1946
rect -3791 -1874 -3757 1946
rect -2533 -1874 -2499 1946
rect -1275 -1874 -1241 1946
rect -17 -1874 17 1946
rect 1241 -1874 1275 1946
rect 2499 -1874 2533 1946
rect 3757 -1874 3791 1946
rect 5015 -1874 5049 1946
rect 6273 -1874 6307 1946
rect 7531 -1874 7565 1946
rect 8789 -1874 8823 1946
rect 10047 -1874 10081 1946
<< mvnsubdiff >>
rect -10227 2584 10227 2596
rect -10227 2550 -8095 2584
rect 8095 2550 10227 2584
rect -10227 2538 10227 2550
rect -10227 -2538 -10169 2538
rect 10169 -2538 10227 2538
rect -10227 -2596 10227 -2538
<< mvnsubdiffcont >>
rect -8095 2550 8095 2584
<< poly >>
rect -10035 2436 -8835 2462
rect -8777 2436 -7577 2462
rect -7519 2436 -6319 2462
rect -6261 2436 -5061 2462
rect -5003 2436 -3803 2462
rect -3745 2436 -2545 2462
rect -2487 2436 -1287 2462
rect -1229 2436 -29 2462
rect 29 2436 1229 2462
rect 1287 2436 2487 2462
rect 2545 2436 3745 2462
rect 3803 2436 5003 2462
rect 5061 2436 6261 2462
rect 6319 2436 7519 2462
rect 7577 2436 8777 2462
rect 8835 2436 10035 2462
rect -10035 -2411 -8835 -2364
rect -10035 -2428 -9961 -2411
rect -9977 -2445 -9961 -2428
rect -8909 -2428 -8835 -2411
rect -8777 -2411 -7577 -2364
rect -8777 -2428 -8703 -2411
rect -8909 -2445 -8893 -2428
rect -9977 -2461 -8893 -2445
rect -8719 -2445 -8703 -2428
rect -7651 -2428 -7577 -2411
rect -7519 -2411 -6319 -2364
rect -7519 -2428 -7445 -2411
rect -7651 -2445 -7635 -2428
rect -8719 -2461 -7635 -2445
rect -7461 -2445 -7445 -2428
rect -6393 -2428 -6319 -2411
rect -6261 -2411 -5061 -2364
rect -6261 -2428 -6187 -2411
rect -6393 -2445 -6377 -2428
rect -7461 -2461 -6377 -2445
rect -6203 -2445 -6187 -2428
rect -5135 -2428 -5061 -2411
rect -5003 -2411 -3803 -2364
rect -5003 -2428 -4929 -2411
rect -5135 -2445 -5119 -2428
rect -6203 -2461 -5119 -2445
rect -4945 -2445 -4929 -2428
rect -3877 -2428 -3803 -2411
rect -3745 -2411 -2545 -2364
rect -3745 -2428 -3671 -2411
rect -3877 -2445 -3861 -2428
rect -4945 -2461 -3861 -2445
rect -3687 -2445 -3671 -2428
rect -2619 -2428 -2545 -2411
rect -2487 -2411 -1287 -2364
rect -2487 -2428 -2413 -2411
rect -2619 -2445 -2603 -2428
rect -3687 -2461 -2603 -2445
rect -2429 -2445 -2413 -2428
rect -1361 -2428 -1287 -2411
rect -1229 -2411 -29 -2364
rect -1229 -2428 -1155 -2411
rect -1361 -2445 -1345 -2428
rect -2429 -2461 -1345 -2445
rect -1171 -2445 -1155 -2428
rect -103 -2428 -29 -2411
rect 29 -2411 1229 -2364
rect 29 -2428 103 -2411
rect -103 -2445 -87 -2428
rect -1171 -2461 -87 -2445
rect 87 -2445 103 -2428
rect 1155 -2428 1229 -2411
rect 1287 -2411 2487 -2364
rect 1287 -2428 1361 -2411
rect 1155 -2445 1171 -2428
rect 87 -2461 1171 -2445
rect 1345 -2445 1361 -2428
rect 2413 -2428 2487 -2411
rect 2545 -2411 3745 -2364
rect 2545 -2428 2619 -2411
rect 2413 -2445 2429 -2428
rect 1345 -2461 2429 -2445
rect 2603 -2445 2619 -2428
rect 3671 -2428 3745 -2411
rect 3803 -2411 5003 -2364
rect 3803 -2428 3877 -2411
rect 3671 -2445 3687 -2428
rect 2603 -2461 3687 -2445
rect 3861 -2445 3877 -2428
rect 4929 -2428 5003 -2411
rect 5061 -2411 6261 -2364
rect 5061 -2428 5135 -2411
rect 4929 -2445 4945 -2428
rect 3861 -2461 4945 -2445
rect 5119 -2445 5135 -2428
rect 6187 -2428 6261 -2411
rect 6319 -2411 7519 -2364
rect 6319 -2428 6393 -2411
rect 6187 -2445 6203 -2428
rect 5119 -2461 6203 -2445
rect 6377 -2445 6393 -2428
rect 7445 -2428 7519 -2411
rect 7577 -2411 8777 -2364
rect 7577 -2428 7651 -2411
rect 7445 -2445 7461 -2428
rect 6377 -2461 7461 -2445
rect 7635 -2445 7651 -2428
rect 8703 -2428 8777 -2411
rect 8835 -2411 10035 -2364
rect 8835 -2428 8909 -2411
rect 8703 -2445 8719 -2428
rect 7635 -2461 8719 -2445
rect 8893 -2445 8909 -2428
rect 9961 -2428 10035 -2411
rect 9961 -2445 9977 -2428
rect 8893 -2461 9977 -2445
<< polycont >>
rect -9961 -2445 -8909 -2411
rect -8703 -2445 -7651 -2411
rect -7445 -2445 -6393 -2411
rect -6187 -2445 -5135 -2411
rect -4929 -2445 -3877 -2411
rect -3671 -2445 -2619 -2411
rect -2413 -2445 -1361 -2411
rect -1155 -2445 -103 -2411
rect 103 -2445 1155 -2411
rect 1361 -2445 2413 -2411
rect 2619 -2445 3671 -2411
rect 3877 -2445 4929 -2411
rect 5135 -2445 6187 -2411
rect 6393 -2445 7445 -2411
rect 7651 -2445 8703 -2411
rect 8909 -2445 9961 -2411
<< locali >>
rect -10215 2550 -8095 2584
rect 8095 2550 10215 2584
rect -10215 -2550 -10181 2550
rect -10081 1946 -10047 1962
rect -10081 -1890 -10047 -1874
rect -8823 1946 -8789 1962
rect -8823 -1890 -8789 -1874
rect -7565 1946 -7531 1962
rect -7565 -1890 -7531 -1874
rect -6307 1946 -6273 1962
rect -6307 -1890 -6273 -1874
rect -5049 1946 -5015 1962
rect -5049 -1890 -5015 -1874
rect -3791 1946 -3757 1962
rect -3791 -1890 -3757 -1874
rect -2533 1946 -2499 1962
rect -2533 -1890 -2499 -1874
rect -1275 1946 -1241 1962
rect -1275 -1890 -1241 -1874
rect -17 1946 17 1962
rect -17 -1890 17 -1874
rect 1241 1946 1275 1962
rect 1241 -1890 1275 -1874
rect 2499 1946 2533 1962
rect 2499 -1890 2533 -1874
rect 3757 1946 3791 1962
rect 3757 -1890 3791 -1874
rect 5015 1946 5049 1962
rect 5015 -1890 5049 -1874
rect 6273 1946 6307 1962
rect 6273 -1890 6307 -1874
rect 7531 1946 7565 1962
rect 7531 -1890 7565 -1874
rect 8789 1946 8823 1962
rect 8789 -1890 8823 -1874
rect 10047 1946 10081 1962
rect 10047 -1890 10081 -1874
rect -9977 -2445 -9961 -2411
rect -8909 -2445 -8893 -2411
rect -8719 -2445 -8703 -2411
rect -7651 -2445 -7635 -2411
rect -7461 -2445 -7445 -2411
rect -6393 -2445 -6377 -2411
rect -6203 -2445 -6187 -2411
rect -5135 -2445 -5119 -2411
rect -4945 -2445 -4929 -2411
rect -3877 -2445 -3861 -2411
rect -3687 -2445 -3671 -2411
rect -2619 -2445 -2603 -2411
rect -2429 -2445 -2413 -2411
rect -1361 -2445 -1345 -2411
rect -1171 -2445 -1155 -2411
rect -103 -2445 -87 -2411
rect 87 -2445 103 -2411
rect 1155 -2445 1171 -2411
rect 1345 -2445 1361 -2411
rect 2413 -2445 2429 -2411
rect 2603 -2445 2619 -2411
rect 3671 -2445 3687 -2411
rect 3861 -2445 3877 -2411
rect 4929 -2445 4945 -2411
rect 5119 -2445 5135 -2411
rect 6187 -2445 6203 -2411
rect 6377 -2445 6393 -2411
rect 7445 -2445 7461 -2411
rect 7635 -2445 7651 -2411
rect 8703 -2445 8719 -2411
rect 8893 -2445 8909 -2411
rect 9961 -2445 9977 -2411
rect 10181 -2550 10215 2550
rect -10215 -2584 10215 -2550
<< viali >>
rect -10081 -1874 -10047 1946
rect -8823 -1874 -8789 1946
rect -7565 -1874 -7531 1946
rect -6307 -1874 -6273 1946
rect -5049 -1874 -5015 1946
rect -3791 -1874 -3757 1946
rect -2533 -1874 -2499 1946
rect -1275 -1874 -1241 1946
rect -17 -1874 17 1946
rect 1241 -1874 1275 1946
rect 2499 -1874 2533 1946
rect 3757 -1874 3791 1946
rect 5015 -1874 5049 1946
rect 6273 -1874 6307 1946
rect 7531 -1874 7565 1946
rect 8789 -1874 8823 1946
rect 10047 -1874 10081 1946
rect -9961 -2445 -8909 -2411
rect -8703 -2445 -7651 -2411
rect -7445 -2445 -6393 -2411
rect -6187 -2445 -5135 -2411
rect -4929 -2445 -3877 -2411
rect -3671 -2445 -2619 -2411
rect -2413 -2445 -1361 -2411
rect -1155 -2445 -103 -2411
rect 103 -2445 1155 -2411
rect 1361 -2445 2413 -2411
rect 2619 -2445 3671 -2411
rect 3877 -2445 4929 -2411
rect 5135 -2445 6187 -2411
rect 6393 -2445 7445 -2411
rect 7651 -2445 8703 -2411
rect 8909 -2445 9961 -2411
<< metal1 >>
rect -10087 1946 -10041 1958
rect -10087 -1874 -10081 1946
rect -10047 -1874 -10041 1946
rect -10087 -1886 -10041 -1874
rect -8829 1946 -8783 1958
rect -8829 -1874 -8823 1946
rect -8789 -1874 -8783 1946
rect -8829 -1886 -8783 -1874
rect -7571 1946 -7525 1958
rect -7571 -1874 -7565 1946
rect -7531 -1874 -7525 1946
rect -7571 -1886 -7525 -1874
rect -6313 1946 -6267 1958
rect -6313 -1874 -6307 1946
rect -6273 -1874 -6267 1946
rect -6313 -1886 -6267 -1874
rect -5055 1946 -5009 1958
rect -5055 -1874 -5049 1946
rect -5015 -1874 -5009 1946
rect -5055 -1886 -5009 -1874
rect -3797 1946 -3751 1958
rect -3797 -1874 -3791 1946
rect -3757 -1874 -3751 1946
rect -3797 -1886 -3751 -1874
rect -2539 1946 -2493 1958
rect -2539 -1874 -2533 1946
rect -2499 -1874 -2493 1946
rect -2539 -1886 -2493 -1874
rect -1281 1946 -1235 1958
rect -1281 -1874 -1275 1946
rect -1241 -1874 -1235 1946
rect -1281 -1886 -1235 -1874
rect -23 1946 23 1958
rect -23 -1874 -17 1946
rect 17 -1874 23 1946
rect -23 -1886 23 -1874
rect 1235 1946 1281 1958
rect 1235 -1874 1241 1946
rect 1275 -1874 1281 1946
rect 1235 -1886 1281 -1874
rect 2493 1946 2539 1958
rect 2493 -1874 2499 1946
rect 2533 -1874 2539 1946
rect 2493 -1886 2539 -1874
rect 3751 1946 3797 1958
rect 3751 -1874 3757 1946
rect 3791 -1874 3797 1946
rect 3751 -1886 3797 -1874
rect 5009 1946 5055 1958
rect 5009 -1874 5015 1946
rect 5049 -1874 5055 1946
rect 5009 -1886 5055 -1874
rect 6267 1946 6313 1958
rect 6267 -1874 6273 1946
rect 6307 -1874 6313 1946
rect 6267 -1886 6313 -1874
rect 7525 1946 7571 1958
rect 7525 -1874 7531 1946
rect 7565 -1874 7571 1946
rect 7525 -1886 7571 -1874
rect 8783 1946 8829 1958
rect 8783 -1874 8789 1946
rect 8823 -1874 8829 1946
rect 8783 -1886 8829 -1874
rect 10041 1946 10087 1958
rect 10041 -1874 10047 1946
rect 10081 -1874 10087 1946
rect 10041 -1886 10087 -1874
rect -9973 -2411 -8897 -2405
rect -9973 -2445 -9961 -2411
rect -8909 -2445 -8897 -2411
rect -9973 -2451 -8897 -2445
rect -8715 -2411 -7639 -2405
rect -8715 -2445 -8703 -2411
rect -7651 -2445 -7639 -2411
rect -8715 -2451 -7639 -2445
rect -7457 -2411 -6381 -2405
rect -7457 -2445 -7445 -2411
rect -6393 -2445 -6381 -2411
rect -7457 -2451 -6381 -2445
rect -6199 -2411 -5123 -2405
rect -6199 -2445 -6187 -2411
rect -5135 -2445 -5123 -2411
rect -6199 -2451 -5123 -2445
rect -4941 -2411 -3865 -2405
rect -4941 -2445 -4929 -2411
rect -3877 -2445 -3865 -2411
rect -4941 -2451 -3865 -2445
rect -3683 -2411 -2607 -2405
rect -3683 -2445 -3671 -2411
rect -2619 -2445 -2607 -2411
rect -3683 -2451 -2607 -2445
rect -2425 -2411 -1349 -2405
rect -2425 -2445 -2413 -2411
rect -1361 -2445 -1349 -2411
rect -2425 -2451 -1349 -2445
rect -1167 -2411 -91 -2405
rect -1167 -2445 -1155 -2411
rect -103 -2445 -91 -2411
rect -1167 -2451 -91 -2445
rect 91 -2411 1167 -2405
rect 91 -2445 103 -2411
rect 1155 -2445 1167 -2411
rect 91 -2451 1167 -2445
rect 1349 -2411 2425 -2405
rect 1349 -2445 1361 -2411
rect 2413 -2445 2425 -2411
rect 1349 -2451 2425 -2445
rect 2607 -2411 3683 -2405
rect 2607 -2445 2619 -2411
rect 3671 -2445 3683 -2411
rect 2607 -2451 3683 -2445
rect 3865 -2411 4941 -2405
rect 3865 -2445 3877 -2411
rect 4929 -2445 4941 -2411
rect 3865 -2451 4941 -2445
rect 5123 -2411 6199 -2405
rect 5123 -2445 5135 -2411
rect 6187 -2445 6199 -2411
rect 5123 -2451 6199 -2445
rect 6381 -2411 7457 -2405
rect 6381 -2445 6393 -2411
rect 7445 -2445 7457 -2411
rect 6381 -2451 7457 -2445
rect 7639 -2411 8715 -2405
rect 7639 -2445 7651 -2411
rect 8703 -2445 8715 -2411
rect 7639 -2451 8715 -2445
rect 8897 -2411 9973 -2405
rect 8897 -2445 8909 -2411
rect 9961 -2445 9973 -2411
rect 8897 -2451 9973 -2445
<< properties >>
string FIXED_BBOX -10198 -2567 10198 2567
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 24.0 l 6.0 m 1 nf 16 diffcov 80 polycov 90 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 80 rlcov 80 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 80 viadrn 80 viagate 90 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
