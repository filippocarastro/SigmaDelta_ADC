magic
tech sky130B
magscale 1 2
timestamp 1666302226
<< nwell >>
rect -858 -10251 858 10251
<< mvpmos >>
rect -600 5154 600 9954
rect -600 118 600 4918
rect -600 -4918 600 -118
rect -600 -9954 600 -5154
<< mvpdiff >>
rect -658 9942 -600 9954
rect -658 5166 -646 9942
rect -612 5166 -600 9942
rect -658 5154 -600 5166
rect 600 9942 658 9954
rect 600 5166 612 9942
rect 646 5166 658 9942
rect 600 5154 658 5166
rect -658 4906 -600 4918
rect -658 130 -646 4906
rect -612 130 -600 4906
rect -658 118 -600 130
rect 600 4906 658 4918
rect 600 130 612 4906
rect 646 130 658 4906
rect 600 118 658 130
rect -658 -130 -600 -118
rect -658 -4906 -646 -130
rect -612 -4906 -600 -130
rect -658 -4918 -600 -4906
rect 600 -130 658 -118
rect 600 -4906 612 -130
rect 646 -4906 658 -130
rect 600 -4918 658 -4906
rect -658 -5166 -600 -5154
rect -658 -9942 -646 -5166
rect -612 -9942 -600 -5166
rect -658 -9954 -600 -9942
rect 600 -5166 658 -5154
rect 600 -9942 612 -5166
rect 646 -9942 658 -5166
rect 600 -9954 658 -9942
<< mvpdiffc >>
rect -646 5166 -612 9942
rect 612 5166 646 9942
rect -646 130 -612 4906
rect 612 130 646 4906
rect -646 -4906 -612 -130
rect 612 -4906 646 -130
rect -646 -9942 -612 -5166
rect 612 -9942 646 -5166
<< mvnsubdiff >>
rect -792 10173 792 10185
rect -792 10139 -684 10173
rect 684 10139 792 10173
rect -792 10127 792 10139
rect -792 10077 -734 10127
rect -792 -10077 -780 10077
rect -746 -10077 -734 10077
rect 734 10077 792 10127
rect -792 -10127 -734 -10077
rect 734 -10077 746 10077
rect 780 -10077 792 10077
rect 734 -10127 792 -10077
rect -792 -10139 792 -10127
rect -792 -10173 -684 -10139
rect 684 -10173 792 -10139
rect -792 -10185 792 -10173
<< mvnsubdiffcont >>
rect -684 10139 684 10173
rect -780 -10077 -746 10077
rect 746 -10077 780 10077
rect -684 -10173 684 -10139
<< poly >>
rect -600 10035 600 10051
rect -600 10001 -584 10035
rect 584 10001 600 10035
rect -600 9954 600 10001
rect -600 5107 600 5154
rect -600 5073 -584 5107
rect 584 5073 600 5107
rect -600 5057 600 5073
rect -600 4999 600 5015
rect -600 4965 -584 4999
rect 584 4965 600 4999
rect -600 4918 600 4965
rect -600 71 600 118
rect -600 37 -584 71
rect 584 37 600 71
rect -600 21 600 37
rect -600 -37 600 -21
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -600 -118 600 -71
rect -600 -4965 600 -4918
rect -600 -4999 -584 -4965
rect 584 -4999 600 -4965
rect -600 -5015 600 -4999
rect -600 -5073 600 -5057
rect -600 -5107 -584 -5073
rect 584 -5107 600 -5073
rect -600 -5154 600 -5107
rect -600 -10001 600 -9954
rect -600 -10035 -584 -10001
rect 584 -10035 600 -10001
rect -600 -10051 600 -10035
<< polycont >>
rect -584 10001 584 10035
rect -584 5073 584 5107
rect -584 4965 584 4999
rect -584 37 584 71
rect -584 -71 584 -37
rect -584 -4999 584 -4965
rect -584 -5107 584 -5073
rect -584 -10035 584 -10001
<< locali >>
rect -780 10139 -684 10173
rect 684 10139 780 10173
rect -780 10077 -746 10139
rect 746 10077 780 10139
rect -600 10001 -584 10035
rect 584 10001 600 10035
rect -646 9942 -612 9958
rect -646 5150 -612 5166
rect 612 9942 646 9958
rect 612 5150 646 5166
rect -600 5073 -584 5107
rect 584 5073 600 5107
rect -600 4965 -584 4999
rect 584 4965 600 4999
rect -646 4906 -612 4922
rect -646 114 -612 130
rect 612 4906 646 4922
rect 612 114 646 130
rect -600 37 -584 71
rect 584 37 600 71
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -646 -130 -612 -114
rect -646 -4922 -612 -4906
rect 612 -130 646 -114
rect 612 -4922 646 -4906
rect -600 -4999 -584 -4965
rect 584 -4999 600 -4965
rect -600 -5107 -584 -5073
rect 584 -5107 600 -5073
rect -646 -5166 -612 -5150
rect -646 -9958 -612 -9942
rect 612 -5166 646 -5150
rect 612 -9958 646 -9942
rect -600 -10035 -584 -10001
rect 584 -10035 600 -10001
rect -780 -10139 -746 -10077
rect 746 -10139 780 -10077
rect -780 -10173 -684 -10139
rect 684 -10173 780 -10139
<< viali >>
rect -584 10001 584 10035
rect -646 5166 -612 9942
rect 612 5166 646 9942
rect -584 5073 584 5107
rect -584 4965 584 4999
rect -646 130 -612 4906
rect 612 130 646 4906
rect -584 37 584 71
rect -584 -71 584 -37
rect -646 -4906 -612 -130
rect 612 -4906 646 -130
rect -584 -4999 584 -4965
rect -584 -5107 584 -5073
rect -646 -9942 -612 -5166
rect 612 -9942 646 -5166
rect -584 -10035 584 -10001
<< metal1 >>
rect -596 10035 596 10041
rect -596 10001 -584 10035
rect 584 10001 596 10035
rect -596 9995 596 10001
rect -652 9942 -606 9954
rect -652 5166 -646 9942
rect -612 5166 -606 9942
rect -652 5154 -606 5166
rect 606 9942 652 9954
rect 606 5166 612 9942
rect 646 5166 652 9942
rect 606 5154 652 5166
rect -596 5107 596 5113
rect -596 5073 -584 5107
rect 584 5073 596 5107
rect -596 5067 596 5073
rect -596 4999 596 5005
rect -596 4965 -584 4999
rect 584 4965 596 4999
rect -596 4959 596 4965
rect -652 4906 -606 4918
rect -652 130 -646 4906
rect -612 130 -606 4906
rect -652 118 -606 130
rect 606 4906 652 4918
rect 606 130 612 4906
rect 646 130 652 4906
rect 606 118 652 130
rect -596 71 596 77
rect -596 37 -584 71
rect 584 37 596 71
rect -596 31 596 37
rect -596 -37 596 -31
rect -596 -71 -584 -37
rect 584 -71 596 -37
rect -596 -77 596 -71
rect -652 -130 -606 -118
rect -652 -4906 -646 -130
rect -612 -4906 -606 -130
rect -652 -4918 -606 -4906
rect 606 -130 652 -118
rect 606 -4906 612 -130
rect 646 -4906 652 -130
rect 606 -4918 652 -4906
rect -596 -4965 596 -4959
rect -596 -4999 -584 -4965
rect 584 -4999 596 -4965
rect -596 -5005 596 -4999
rect -596 -5073 596 -5067
rect -596 -5107 -584 -5073
rect 584 -5107 596 -5073
rect -596 -5113 596 -5107
rect -652 -5166 -606 -5154
rect -652 -9942 -646 -5166
rect -612 -9942 -606 -5166
rect -652 -9954 -606 -9942
rect 606 -5166 652 -5154
rect 606 -9942 612 -5166
rect 646 -9942 652 -5166
rect 606 -9954 652 -9942
rect -596 -10001 596 -9995
rect -596 -10035 -584 -10001
rect 584 -10035 596 -10001
rect -596 -10041 596 -10035
<< properties >>
string FIXED_BBOX -763 -10156 763 10156
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 24.0 l 6.0 m 4 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
