magic
tech sky130B
magscale 1 2
timestamp 1667120857
<< nwell >>
rect -2745 -2662 2745 2662
<< mvpmos >>
rect -2487 -2436 -1287 2364
rect -1229 -2436 -29 2364
rect 29 -2436 1229 2364
rect 1287 -2436 2487 2364
<< mvpdiff >>
rect -2545 2352 -2487 2364
rect -2545 -2424 -2533 2352
rect -2499 -2424 -2487 2352
rect -2545 -2436 -2487 -2424
rect -1287 2352 -1229 2364
rect -1287 -2424 -1275 2352
rect -1241 -2424 -1229 2352
rect -1287 -2436 -1229 -2424
rect -29 2352 29 2364
rect -29 -2424 -17 2352
rect 17 -2424 29 2352
rect -29 -2436 29 -2424
rect 1229 2352 1287 2364
rect 1229 -2424 1241 2352
rect 1275 -2424 1287 2352
rect 1229 -2436 1287 -2424
rect 2487 2352 2545 2364
rect 2487 -2424 2499 2352
rect 2533 -2424 2545 2352
rect 2487 -2436 2545 -2424
<< mvpdiffc >>
rect -2533 -2424 -2499 2352
rect -1275 -2424 -1241 2352
rect -17 -2424 17 2352
rect 1241 -2424 1275 2352
rect 2499 -2424 2533 2352
<< mvnsubdiff >>
rect -2679 2584 2679 2596
rect -2679 2550 -2571 2584
rect 2571 2550 2679 2584
rect -2679 2538 2679 2550
rect -2679 2488 -2621 2538
rect -2679 -2488 -2667 2488
rect -2633 -2488 -2621 2488
rect 2621 2488 2679 2538
rect -2679 -2538 -2621 -2488
rect 2621 -2488 2633 2488
rect 2667 -2488 2679 2488
rect 2621 -2538 2679 -2488
rect -2679 -2550 2679 -2538
rect -2679 -2584 -2571 -2550
rect 2571 -2584 2679 -2550
rect -2679 -2596 2679 -2584
<< mvnsubdiffcont >>
rect -2571 2550 2571 2584
rect -2667 -2488 -2633 2488
rect 2633 -2488 2667 2488
rect -2571 -2584 2571 -2550
<< poly >>
rect -2487 2445 -1287 2461
rect -2487 2411 -2471 2445
rect -1303 2411 -1287 2445
rect -2487 2364 -1287 2411
rect -1229 2445 -29 2461
rect -1229 2411 -1213 2445
rect -45 2411 -29 2445
rect -1229 2364 -29 2411
rect 29 2445 1229 2461
rect 29 2411 45 2445
rect 1213 2411 1229 2445
rect 29 2364 1229 2411
rect 1287 2445 2487 2461
rect 1287 2411 1303 2445
rect 2471 2411 2487 2445
rect 1287 2364 2487 2411
rect -2487 -2462 -1287 -2436
rect -1229 -2462 -29 -2436
rect 29 -2462 1229 -2436
rect 1287 -2462 2487 -2436
<< polycont >>
rect -2471 2411 -1303 2445
rect -1213 2411 -45 2445
rect 45 2411 1213 2445
rect 1303 2411 2471 2445
<< locali >>
rect -2667 2550 -2571 2584
rect 2571 2550 2667 2584
rect -2667 2488 -2633 2550
rect 2633 2488 2667 2550
rect -2487 2411 -2471 2445
rect -1303 2411 -1287 2445
rect -1229 2411 -1213 2445
rect -45 2411 -29 2445
rect 29 2411 45 2445
rect 1213 2411 1229 2445
rect 1287 2411 1303 2445
rect 2471 2411 2487 2445
rect -2533 2352 -2499 2368
rect -2533 -2440 -2499 -2424
rect -1275 2352 -1241 2368
rect -1275 -2440 -1241 -2424
rect -17 2352 17 2368
rect -17 -2440 17 -2424
rect 1241 2352 1275 2368
rect 1241 -2440 1275 -2424
rect 2499 2352 2533 2368
rect 2499 -2440 2533 -2424
rect -2667 -2550 -2633 -2488
rect 2633 -2550 2667 -2488
rect -2667 -2584 -2571 -2550
rect 2571 -2584 2667 -2550
<< viali >>
rect -2471 2411 -1303 2445
rect -1213 2411 -45 2445
rect 45 2411 1213 2445
rect 1303 2411 2471 2445
rect -2533 -2424 -2499 2352
rect -1275 -2424 -1241 2352
rect -17 -2424 17 2352
rect 1241 -2424 1275 2352
rect 2499 -2424 2533 2352
<< metal1 >>
rect -2483 2445 -1291 2451
rect -2483 2411 -2471 2445
rect -1303 2411 -1291 2445
rect -2483 2405 -1291 2411
rect -1225 2445 -33 2451
rect -1225 2411 -1213 2445
rect -45 2411 -33 2445
rect -1225 2405 -33 2411
rect 33 2445 1225 2451
rect 33 2411 45 2445
rect 1213 2411 1225 2445
rect 33 2405 1225 2411
rect 1291 2445 2483 2451
rect 1291 2411 1303 2445
rect 2471 2411 2483 2445
rect 1291 2405 2483 2411
rect -2539 2352 -2493 2364
rect -2539 -2424 -2533 2352
rect -2499 -2424 -2493 2352
rect -2539 -2436 -2493 -2424
rect -1281 2352 -1235 2364
rect -1281 -2424 -1275 2352
rect -1241 -2424 -1235 2352
rect -1281 -2436 -1235 -2424
rect -23 2352 23 2364
rect -23 -2424 -17 2352
rect 17 -2424 23 2352
rect -23 -2436 23 -2424
rect 1235 2352 1281 2364
rect 1235 -2424 1241 2352
rect 1275 -2424 1281 2352
rect 1235 -2436 1281 -2424
rect 2493 2352 2539 2364
rect 2493 -2424 2499 2352
rect 2533 -2424 2539 2352
rect 2493 -2436 2539 -2424
<< properties >>
string FIXED_BBOX -2650 -2567 2650 2567
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 24.0 l 6.0 m 1 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
