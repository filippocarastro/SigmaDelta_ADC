magic
tech sky130B
timestamp 1667069721
<< pwell >>
rect -1672 -2529 1672 2529
<< mvnmos >>
rect -1558 -2400 -958 2400
rect -929 -2400 -329 2400
rect -300 -2400 300 2400
rect 329 -2400 929 2400
rect 958 -2400 1558 2400
<< mvndiff >>
rect -1587 2394 -1558 2400
rect -1587 -2394 -1581 2394
rect -1564 -2394 -1558 2394
rect -1587 -2400 -1558 -2394
rect -958 2394 -929 2400
rect -958 -2394 -952 2394
rect -935 -2394 -929 2394
rect -958 -2400 -929 -2394
rect -329 2394 -300 2400
rect -329 -2394 -323 2394
rect -306 -2394 -300 2394
rect -329 -2400 -300 -2394
rect 300 2394 329 2400
rect 300 -2394 306 2394
rect 323 -2394 329 2394
rect 300 -2400 329 -2394
rect 929 2394 958 2400
rect 929 -2394 935 2394
rect 952 -2394 958 2394
rect 929 -2400 958 -2394
rect 1558 2394 1587 2400
rect 1558 -2394 1564 2394
rect 1581 -2394 1587 2394
rect 1558 -2400 1587 -2394
<< mvndiffc >>
rect -1581 -2394 -1564 2394
rect -952 -2394 -935 2394
rect -323 -2394 -306 2394
rect 306 -2394 323 2394
rect 935 -2394 952 2394
rect 1564 -2394 1581 2394
<< mvpsubdiff >>
rect -1654 2505 1654 2511
rect -1654 2488 -1600 2505
rect 1600 2488 1654 2505
rect -1654 2482 1654 2488
rect -1654 2457 -1625 2482
rect -1654 -2457 -1648 2457
rect -1631 -2457 -1625 2457
rect 1625 2457 1654 2482
rect -1654 -2482 -1625 -2457
rect 1625 -2457 1631 2457
rect 1648 -2457 1654 2457
rect 1625 -2482 1654 -2457
rect -1654 -2488 1654 -2482
rect -1654 -2505 -1600 -2488
rect 1600 -2505 1654 -2488
rect -1654 -2511 1654 -2505
<< mvpsubdiffcont >>
rect -1600 2488 1600 2505
rect -1648 -2457 -1631 2457
rect 1631 -2457 1648 2457
rect -1600 -2505 1600 -2488
<< poly >>
rect -1558 2436 -958 2444
rect -1558 2419 -1550 2436
rect -966 2419 -958 2436
rect -1558 2400 -958 2419
rect -929 2436 -329 2444
rect -929 2419 -921 2436
rect -337 2419 -329 2436
rect -929 2400 -329 2419
rect -300 2436 300 2444
rect -300 2419 -292 2436
rect 292 2419 300 2436
rect -300 2400 300 2419
rect 329 2436 929 2444
rect 329 2419 337 2436
rect 921 2419 929 2436
rect 329 2400 929 2419
rect 958 2436 1558 2444
rect 958 2419 966 2436
rect 1550 2419 1558 2436
rect 958 2400 1558 2419
rect -1558 -2419 -958 -2400
rect -1558 -2436 -1550 -2419
rect -966 -2436 -958 -2419
rect -1558 -2444 -958 -2436
rect -929 -2419 -329 -2400
rect -929 -2436 -921 -2419
rect -337 -2436 -329 -2419
rect -929 -2444 -329 -2436
rect -300 -2419 300 -2400
rect -300 -2436 -292 -2419
rect 292 -2436 300 -2419
rect -300 -2444 300 -2436
rect 329 -2419 929 -2400
rect 329 -2436 337 -2419
rect 921 -2436 929 -2419
rect 329 -2444 929 -2436
rect 958 -2419 1558 -2400
rect 958 -2436 966 -2419
rect 1550 -2436 1558 -2419
rect 958 -2444 1558 -2436
<< polycont >>
rect -1550 2419 -966 2436
rect -921 2419 -337 2436
rect -292 2419 292 2436
rect 337 2419 921 2436
rect 966 2419 1550 2436
rect -1550 -2436 -966 -2419
rect -921 -2436 -337 -2419
rect -292 -2436 292 -2419
rect 337 -2436 921 -2419
rect 966 -2436 1550 -2419
<< locali >>
rect -1648 2488 -1600 2505
rect 1600 2488 1648 2505
rect -1648 2457 -1631 2488
rect 1631 2457 1648 2488
rect -1558 2419 -1550 2436
rect -966 2419 -958 2436
rect -929 2419 -921 2436
rect -337 2419 -329 2436
rect -300 2419 -292 2436
rect 292 2419 300 2436
rect 329 2419 337 2436
rect 921 2419 929 2436
rect 958 2419 966 2436
rect 1550 2419 1558 2436
rect -1581 2394 -1564 2402
rect -1581 -2402 -1564 -2394
rect -952 2394 -935 2402
rect -952 -2402 -935 -2394
rect -323 2394 -306 2402
rect -323 -2402 -306 -2394
rect 306 2394 323 2402
rect 306 -2402 323 -2394
rect 935 2394 952 2402
rect 935 -2402 952 -2394
rect 1564 2394 1581 2402
rect 1564 -2402 1581 -2394
rect -1558 -2436 -1550 -2419
rect -966 -2436 -958 -2419
rect -929 -2436 -921 -2419
rect -337 -2436 -329 -2419
rect -300 -2436 -292 -2419
rect 292 -2436 300 -2419
rect 329 -2436 337 -2419
rect 921 -2436 929 -2419
rect 958 -2436 966 -2419
rect 1550 -2436 1558 -2419
rect -1648 -2488 -1631 -2457
rect 1631 -2488 1648 -2457
rect -1648 -2505 -1600 -2488
rect 1600 -2505 1648 -2488
<< viali >>
rect -1550 2419 -966 2436
rect -921 2419 -337 2436
rect -292 2419 292 2436
rect 337 2419 921 2436
rect 966 2419 1550 2436
rect -1581 -2394 -1564 2394
rect -952 -2394 -935 2394
rect -323 -2394 -306 2394
rect 306 -2394 323 2394
rect 935 -2394 952 2394
rect 1564 -2394 1581 2394
rect -1550 -2436 -966 -2419
rect -921 -2436 -337 -2419
rect -292 -2436 292 -2419
rect 337 -2436 921 -2419
rect 966 -2436 1550 -2419
<< metal1 >>
rect -1556 2436 -960 2439
rect -1556 2419 -1550 2436
rect -966 2419 -960 2436
rect -1556 2416 -960 2419
rect -927 2436 -331 2439
rect -927 2419 -921 2436
rect -337 2419 -331 2436
rect -927 2416 -331 2419
rect -298 2436 298 2439
rect -298 2419 -292 2436
rect 292 2419 298 2436
rect -298 2416 298 2419
rect 331 2436 927 2439
rect 331 2419 337 2436
rect 921 2419 927 2436
rect 331 2416 927 2419
rect 960 2436 1556 2439
rect 960 2419 966 2436
rect 1550 2419 1556 2436
rect 960 2416 1556 2419
rect -1584 2394 -1561 2400
rect -1584 -2394 -1581 2394
rect -1564 -2394 -1561 2394
rect -1584 -2400 -1561 -2394
rect -955 2394 -932 2400
rect -955 -2394 -952 2394
rect -935 -2394 -932 2394
rect -955 -2400 -932 -2394
rect -326 2394 -303 2400
rect -326 -2394 -323 2394
rect -306 -2394 -303 2394
rect -326 -2400 -303 -2394
rect 303 2394 326 2400
rect 303 -2394 306 2394
rect 323 -2394 326 2394
rect 303 -2400 326 -2394
rect 932 2394 955 2400
rect 932 -2394 935 2394
rect 952 -2394 955 2394
rect 932 -2400 955 -2394
rect 1561 2394 1584 2400
rect 1561 -2394 1564 2394
rect 1581 -2394 1584 2394
rect 1561 -2400 1584 -2394
rect -1556 -2419 -960 -2416
rect -1556 -2436 -1550 -2419
rect -966 -2436 -960 -2419
rect -1556 -2439 -960 -2436
rect -927 -2419 -331 -2416
rect -927 -2436 -921 -2419
rect -337 -2436 -331 -2419
rect -927 -2439 -331 -2436
rect -298 -2419 298 -2416
rect -298 -2436 -292 -2419
rect 292 -2436 298 -2419
rect -298 -2439 298 -2436
rect 331 -2419 927 -2416
rect 331 -2436 337 -2419
rect 921 -2436 927 -2419
rect 331 -2439 927 -2436
rect 960 -2419 1556 -2416
rect 960 -2436 966 -2419
rect 1550 -2436 1556 -2419
rect 960 -2439 1556 -2436
<< properties >>
string FIXED_BBOX -1639 -2496 1639 2496
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 48.0 l 6.0 m 1 nf 5 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
