magic
tech sky130B
magscale 1 2
timestamp 1666302226
<< nwell >>
rect -4003 -3497 4003 3497
<< mvpmos >>
rect -3745 -3200 -2545 3200
rect -2487 -3200 -1287 3200
rect -1229 -3200 -29 3200
rect 29 -3200 1229 3200
rect 1287 -3200 2487 3200
rect 2545 -3200 3745 3200
<< mvpdiff >>
rect -3803 3188 -3745 3200
rect -3803 -3188 -3791 3188
rect -3757 -3188 -3745 3188
rect -3803 -3200 -3745 -3188
rect -2545 3188 -2487 3200
rect -2545 -3188 -2533 3188
rect -2499 -3188 -2487 3188
rect -2545 -3200 -2487 -3188
rect -1287 3188 -1229 3200
rect -1287 -3188 -1275 3188
rect -1241 -3188 -1229 3188
rect -1287 -3200 -1229 -3188
rect -29 3188 29 3200
rect -29 -3188 -17 3188
rect 17 -3188 29 3188
rect -29 -3200 29 -3188
rect 1229 3188 1287 3200
rect 1229 -3188 1241 3188
rect 1275 -3188 1287 3188
rect 1229 -3200 1287 -3188
rect 2487 3188 2545 3200
rect 2487 -3188 2499 3188
rect 2533 -3188 2545 3188
rect 2487 -3200 2545 -3188
rect 3745 3188 3803 3200
rect 3745 -3188 3757 3188
rect 3791 -3188 3803 3188
rect 3745 -3200 3803 -3188
<< mvpdiffc >>
rect -3791 -3188 -3757 3188
rect -2533 -3188 -2499 3188
rect -1275 -3188 -1241 3188
rect -17 -3188 17 3188
rect 1241 -3188 1275 3188
rect 2499 -3188 2533 3188
rect 3757 -3188 3791 3188
<< mvnsubdiff >>
rect -3937 3419 3937 3431
rect -3937 3385 -3829 3419
rect 3829 3385 3937 3419
rect -3937 3373 3937 3385
rect -3937 3323 -3879 3373
rect -3937 -3323 -3925 3323
rect -3891 -3323 -3879 3323
rect 3879 3323 3937 3373
rect -3937 -3373 -3879 -3323
rect 3879 -3323 3891 3323
rect 3925 -3323 3937 3323
rect 3879 -3373 3937 -3323
rect -3937 -3385 3937 -3373
rect -3937 -3419 -3829 -3385
rect 3829 -3419 3937 -3385
rect -3937 -3431 3937 -3419
<< mvnsubdiffcont >>
rect -3829 3385 3829 3419
rect -3925 -3323 -3891 3323
rect 3891 -3323 3925 3323
rect -3829 -3419 3829 -3385
<< poly >>
rect -3745 3281 -2545 3297
rect -3745 3247 -3729 3281
rect -2561 3247 -2545 3281
rect -3745 3200 -2545 3247
rect -2487 3281 -1287 3297
rect -2487 3247 -2471 3281
rect -1303 3247 -1287 3281
rect -2487 3200 -1287 3247
rect -1229 3281 -29 3297
rect -1229 3247 -1213 3281
rect -45 3247 -29 3281
rect -1229 3200 -29 3247
rect 29 3281 1229 3297
rect 29 3247 45 3281
rect 1213 3247 1229 3281
rect 29 3200 1229 3247
rect 1287 3281 2487 3297
rect 1287 3247 1303 3281
rect 2471 3247 2487 3281
rect 1287 3200 2487 3247
rect 2545 3281 3745 3297
rect 2545 3247 2561 3281
rect 3729 3247 3745 3281
rect 2545 3200 3745 3247
rect -3745 -3247 -2545 -3200
rect -3745 -3281 -3729 -3247
rect -2561 -3281 -2545 -3247
rect -3745 -3297 -2545 -3281
rect -2487 -3247 -1287 -3200
rect -2487 -3281 -2471 -3247
rect -1303 -3281 -1287 -3247
rect -2487 -3297 -1287 -3281
rect -1229 -3247 -29 -3200
rect -1229 -3281 -1213 -3247
rect -45 -3281 -29 -3247
rect -1229 -3297 -29 -3281
rect 29 -3247 1229 -3200
rect 29 -3281 45 -3247
rect 1213 -3281 1229 -3247
rect 29 -3297 1229 -3281
rect 1287 -3247 2487 -3200
rect 1287 -3281 1303 -3247
rect 2471 -3281 2487 -3247
rect 1287 -3297 2487 -3281
rect 2545 -3247 3745 -3200
rect 2545 -3281 2561 -3247
rect 3729 -3281 3745 -3247
rect 2545 -3297 3745 -3281
<< polycont >>
rect -3729 3247 -2561 3281
rect -2471 3247 -1303 3281
rect -1213 3247 -45 3281
rect 45 3247 1213 3281
rect 1303 3247 2471 3281
rect 2561 3247 3729 3281
rect -3729 -3281 -2561 -3247
rect -2471 -3281 -1303 -3247
rect -1213 -3281 -45 -3247
rect 45 -3281 1213 -3247
rect 1303 -3281 2471 -3247
rect 2561 -3281 3729 -3247
<< locali >>
rect -3925 3385 -3829 3419
rect 3829 3385 3925 3419
rect -3925 3323 -3891 3385
rect 3891 3323 3925 3385
rect -3745 3247 -3729 3281
rect -2561 3247 -2545 3281
rect -2487 3247 -2471 3281
rect -1303 3247 -1287 3281
rect -1229 3247 -1213 3281
rect -45 3247 -29 3281
rect 29 3247 45 3281
rect 1213 3247 1229 3281
rect 1287 3247 1303 3281
rect 2471 3247 2487 3281
rect 2545 3247 2561 3281
rect 3729 3247 3745 3281
rect -3791 3188 -3757 3204
rect -3791 -3204 -3757 -3188
rect -2533 3188 -2499 3204
rect -2533 -3204 -2499 -3188
rect -1275 3188 -1241 3204
rect -1275 -3204 -1241 -3188
rect -17 3188 17 3204
rect -17 -3204 17 -3188
rect 1241 3188 1275 3204
rect 1241 -3204 1275 -3188
rect 2499 3188 2533 3204
rect 2499 -3204 2533 -3188
rect 3757 3188 3791 3204
rect 3757 -3204 3791 -3188
rect -3745 -3281 -3729 -3247
rect -2561 -3281 -2545 -3247
rect -2487 -3281 -2471 -3247
rect -1303 -3281 -1287 -3247
rect -1229 -3281 -1213 -3247
rect -45 -3281 -29 -3247
rect 29 -3281 45 -3247
rect 1213 -3281 1229 -3247
rect 1287 -3281 1303 -3247
rect 2471 -3281 2487 -3247
rect 2545 -3281 2561 -3247
rect 3729 -3281 3745 -3247
rect -3925 -3385 -3891 -3323
rect 3891 -3385 3925 -3323
rect -3925 -3419 -3829 -3385
rect 3829 -3419 3925 -3385
<< viali >>
rect -3729 3247 -2561 3281
rect -2471 3247 -1303 3281
rect -1213 3247 -45 3281
rect 45 3247 1213 3281
rect 1303 3247 2471 3281
rect 2561 3247 3729 3281
rect -3791 -3188 -3757 3188
rect -2533 -3188 -2499 3188
rect -1275 -3188 -1241 3188
rect -17 -3188 17 3188
rect 1241 -3188 1275 3188
rect 2499 -3188 2533 3188
rect 3757 -3188 3791 3188
rect -3729 -3281 -2561 -3247
rect -2471 -3281 -1303 -3247
rect -1213 -3281 -45 -3247
rect 45 -3281 1213 -3247
rect 1303 -3281 2471 -3247
rect 2561 -3281 3729 -3247
<< metal1 >>
rect -3741 3281 -2549 3287
rect -3741 3247 -3729 3281
rect -2561 3247 -2549 3281
rect -3741 3241 -2549 3247
rect -2483 3281 -1291 3287
rect -2483 3247 -2471 3281
rect -1303 3247 -1291 3281
rect -2483 3241 -1291 3247
rect -1225 3281 -33 3287
rect -1225 3247 -1213 3281
rect -45 3247 -33 3281
rect -1225 3241 -33 3247
rect 33 3281 1225 3287
rect 33 3247 45 3281
rect 1213 3247 1225 3281
rect 33 3241 1225 3247
rect 1291 3281 2483 3287
rect 1291 3247 1303 3281
rect 2471 3247 2483 3281
rect 1291 3241 2483 3247
rect 2549 3281 3741 3287
rect 2549 3247 2561 3281
rect 3729 3247 3741 3281
rect 2549 3241 3741 3247
rect -3797 3188 -3751 3200
rect -3797 -3188 -3791 3188
rect -3757 -3188 -3751 3188
rect -3797 -3200 -3751 -3188
rect -2539 3188 -2493 3200
rect -2539 -3188 -2533 3188
rect -2499 -3188 -2493 3188
rect -2539 -3200 -2493 -3188
rect -1281 3188 -1235 3200
rect -1281 -3188 -1275 3188
rect -1241 -3188 -1235 3188
rect -1281 -3200 -1235 -3188
rect -23 3188 23 3200
rect -23 -3188 -17 3188
rect 17 -3188 23 3188
rect -23 -3200 23 -3188
rect 1235 3188 1281 3200
rect 1235 -3188 1241 3188
rect 1275 -3188 1281 3188
rect 1235 -3200 1281 -3188
rect 2493 3188 2539 3200
rect 2493 -3188 2499 3188
rect 2533 -3188 2539 3188
rect 2493 -3200 2539 -3188
rect 3751 3188 3797 3200
rect 3751 -3188 3757 3188
rect 3791 -3188 3797 3188
rect 3751 -3200 3797 -3188
rect -3741 -3247 -2549 -3241
rect -3741 -3281 -3729 -3247
rect -2561 -3281 -2549 -3247
rect -3741 -3287 -2549 -3281
rect -2483 -3247 -1291 -3241
rect -2483 -3281 -2471 -3247
rect -1303 -3281 -1291 -3247
rect -2483 -3287 -1291 -3281
rect -1225 -3247 -33 -3241
rect -1225 -3281 -1213 -3247
rect -45 -3281 -33 -3247
rect -1225 -3287 -33 -3281
rect 33 -3247 1225 -3241
rect 33 -3281 45 -3247
rect 1213 -3281 1225 -3247
rect 33 -3287 1225 -3281
rect 1291 -3247 2483 -3241
rect 1291 -3281 1303 -3247
rect 2471 -3281 2483 -3247
rect 1291 -3287 2483 -3281
rect 2549 -3247 3741 -3241
rect 2549 -3281 2561 -3247
rect 3729 -3281 3741 -3247
rect 2549 -3287 3741 -3281
<< properties >>
string FIXED_BBOX -3908 -3402 3908 3402
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 6.0 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
