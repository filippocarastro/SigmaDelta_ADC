magic
tech sky130B
magscale 1 2
timestamp 1667415230
<< metal1 >>
rect 11988 35104 44904 36638
rect 11988 35102 42004 35104
rect 42778 35102 44904 35104
rect 13556 34380 13562 34880
rect 14062 34380 15292 34880
rect 14792 30642 15292 34380
rect 35100 30655 35750 35102
rect 36302 34366 36841 34660
rect 36302 31243 36835 34366
rect 35912 30710 35918 31243
rect 36451 30710 36835 31243
rect 41524 30702 42004 35102
rect 42378 34378 42752 34680
rect 14835 30290 37650 30291
rect 42378 30290 42680 34378
rect 43912 30614 44884 35102
rect 14835 30287 43690 30290
rect 14835 30248 43857 30287
rect 14835 29801 43858 30248
rect 14835 29499 45329 29801
rect 14835 29406 43858 29499
rect 14835 29404 43690 29406
rect 36006 29308 36394 29314
rect 13848 28028 14048 28228
rect 26604 28092 34477 28498
rect 36006 27896 36394 28920
rect 36758 28190 45408 28602
rect 14777 25544 24229 25846
rect 20736 25226 21472 25234
rect 13316 16036 14520 24924
rect 19882 24490 20736 24748
rect 19882 24294 21472 24490
rect 23927 24360 24229 25544
rect 23926 24354 24230 24360
rect 19882 23896 21428 24294
rect 21826 23896 21832 24294
rect 23926 24044 24230 24050
rect 19882 16632 21472 23896
rect 27514 21206 28100 27878
rect 34092 22979 36394 27896
rect 34092 22573 36397 22979
rect 27514 20844 43715 21206
rect 27514 16551 28100 20844
rect 28908 16036 29454 20420
rect 41680 16593 42648 20404
rect 43766 16860 44222 27916
rect 41680 16036 42661 16593
rect 43766 16404 44914 16860
rect 45370 16404 45376 16860
rect 43766 16198 44222 16404
rect 11752 16014 43830 16036
rect 11752 13988 45222 16014
<< via1 >>
rect 13562 34380 14062 34880
rect 35918 30710 36451 31243
rect 36006 28920 36394 29308
rect 20736 24490 21472 25226
rect 21428 23896 21826 24294
rect 23926 24050 24230 24354
rect 44914 16404 45370 16860
<< metal2 >>
rect 13560 34880 14297 34994
rect 13560 34380 13562 34880
rect 14062 34380 14297 34880
rect 13560 28435 14297 34380
rect 35918 31243 36451 31249
rect 35918 29308 36451 30710
rect 35918 28920 36006 29308
rect 36394 28920 36451 29308
rect 35918 28910 36451 28920
rect 13560 27698 21473 28435
rect 20736 25226 21472 27698
rect 20730 24490 20736 25226
rect 21472 24490 21478 25226
rect 21428 24294 21826 24300
rect 21826 23896 22053 24294
rect 22451 23896 22460 24294
rect 23920 24050 23926 24354
rect 24230 24050 24236 24354
rect 21428 23890 21826 23896
rect 23926 20950 24230 24050
rect 23742 20550 24230 20950
rect 23742 16860 24198 20550
rect 44914 16860 45370 16866
rect 23742 16404 44914 16860
rect 44914 16398 45370 16404
<< via2 >>
rect 22053 23896 22451 24294
<< metal3 >>
rect 22048 24294 22456 24299
rect 22048 23896 22053 24294
rect 22451 23896 23310 24294
rect 22048 23891 22456 23896
rect 22643 23666 23310 23896
rect 22642 22692 23310 23666
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1667223724
transform 1 0 24090 0 1 20400
box -3150 -3100 3149 3100
use sky130_fd_pr__nfet_g5v0d10v5_U4FG9E  XM1
timestamp 1667224822
transform 1 0 43184 0 1 18477
box -828 -2627 828 2627
use sky130_fd_pr__pfet_g5v0d10v5_VS8EJU  XM2
timestamp 1667224016
transform 1 0 31046 0 -1 25238
box -3374 -3462 3374 3462
use sky130_fd_pr__nfet_01v8_45ERJ4  XM3
timestamp 1667324858
transform 1 0 28674 0 1 18483
box -796 -2579 796 2579
use sky130_fd_pr__pfet_g5v0d10v5_VS8V9Y  XM4
timestamp 1667223724
transform 1 0 40119 0 1 25266
box -4003 -3462 4003 3462
use sky130_fd_pr__pfet_g5v0d10v5_VSGFLU  XM5
timestamp 1667223724
transform -1 0 39185 0 -1 32696
box -2745 -2662 2745 2662
use sky130_fd_pr__pfet_g5v0d10v5_YHBQGB  XM6
timestamp 1667223724
transform 1 0 25251 0 1 32660
box -10293 -2662 10293 2662
use sky130_fd_pr__nfet_g5v0d10v5_8VPWNZ  XM7
timestamp 1667325532
transform 1 0 17202 0 1 20921
box -3344 -5027 3344 5027
use sky130_fd_pr__pfet_g5v0d10v5_VSGNQY  XM8
timestamp 1667223724
transform 1 0 43332 0 1 32694
box -858 -2662 858 2662
<< labels >>
flabel metal1 12642 35948 12842 36148 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 45106 29566 45306 29766 0 FreeSans 256 0 0 0 Ibias
port 4 nsew
flabel metal1 45192 28196 45392 28396 0 FreeSans 256 0 0 0 Vinp
port 1 nsew
flabel metal1 26604 28092 26804 28292 0 FreeSans 256 0 0 0 Vinn
port 0 nsew
flabel metal1 44802 14338 45002 14538 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 13848 28028 14048 28228 0 FreeSans 256 0 0 0 Vout
port 5 nsew
<< end >>
