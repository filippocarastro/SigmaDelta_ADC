magic
tech sky130B
magscale 1 2
timestamp 1667120857
<< nwell >>
rect -2116 -10027 2116 10027
<< mvpmos >>
rect -1858 3329 -658 9729
rect -600 3329 600 9729
rect 658 3329 1858 9729
rect -1858 -3236 -658 3164
rect -600 -3236 600 3164
rect 658 -3236 1858 3164
rect -1858 -9801 -658 -3401
rect -600 -9801 600 -3401
rect 658 -9801 1858 -3401
<< mvpdiff >>
rect -1916 9717 -1858 9729
rect -1916 3341 -1904 9717
rect -1870 3341 -1858 9717
rect -1916 3329 -1858 3341
rect -658 9717 -600 9729
rect -658 3341 -646 9717
rect -612 3341 -600 9717
rect -658 3329 -600 3341
rect 600 9717 658 9729
rect 600 3341 612 9717
rect 646 3341 658 9717
rect 600 3329 658 3341
rect 1858 9717 1916 9729
rect 1858 3341 1870 9717
rect 1904 3341 1916 9717
rect 1858 3329 1916 3341
rect -1916 3152 -1858 3164
rect -1916 -3224 -1904 3152
rect -1870 -3224 -1858 3152
rect -1916 -3236 -1858 -3224
rect -658 3152 -600 3164
rect -658 -3224 -646 3152
rect -612 -3224 -600 3152
rect -658 -3236 -600 -3224
rect 600 3152 658 3164
rect 600 -3224 612 3152
rect 646 -3224 658 3152
rect 600 -3236 658 -3224
rect 1858 3152 1916 3164
rect 1858 -3224 1870 3152
rect 1904 -3224 1916 3152
rect 1858 -3236 1916 -3224
rect -1916 -3413 -1858 -3401
rect -1916 -9789 -1904 -3413
rect -1870 -9789 -1858 -3413
rect -1916 -9801 -1858 -9789
rect -658 -3413 -600 -3401
rect -658 -9789 -646 -3413
rect -612 -9789 -600 -3413
rect -658 -9801 -600 -9789
rect 600 -3413 658 -3401
rect 600 -9789 612 -3413
rect 646 -9789 658 -3413
rect 600 -9801 658 -9789
rect 1858 -3413 1916 -3401
rect 1858 -9789 1870 -3413
rect 1904 -9789 1916 -3413
rect 1858 -9801 1916 -9789
<< mvpdiffc >>
rect -1904 3341 -1870 9717
rect -646 3341 -612 9717
rect 612 3341 646 9717
rect 1870 3341 1904 9717
rect -1904 -3224 -1870 3152
rect -646 -3224 -612 3152
rect 612 -3224 646 3152
rect 1870 -3224 1904 3152
rect -1904 -9789 -1870 -3413
rect -646 -9789 -612 -3413
rect 612 -9789 646 -3413
rect 1870 -9789 1904 -3413
<< mvnsubdiff >>
rect -2050 9949 2050 9961
rect -2050 9915 -1942 9949
rect 1942 9915 2050 9949
rect -2050 9903 2050 9915
rect -2050 9853 -1992 9903
rect -2050 -9853 -2038 9853
rect -2004 -9853 -1992 9853
rect 1992 9853 2050 9903
rect -2050 -9903 -1992 -9853
rect 1992 -9853 2004 9853
rect 2038 -9853 2050 9853
rect 1992 -9903 2050 -9853
rect -2050 -9915 2050 -9903
rect -2050 -9949 -1942 -9915
rect 1942 -9949 2050 -9915
rect -2050 -9961 2050 -9949
<< mvnsubdiffcont >>
rect -1942 9915 1942 9949
rect -2038 -9853 -2004 9853
rect 2004 -9853 2038 9853
rect -1942 -9949 1942 -9915
<< poly >>
rect -1858 9810 -658 9826
rect -1858 9776 -1842 9810
rect -674 9776 -658 9810
rect -1858 9729 -658 9776
rect -600 9810 600 9826
rect -600 9776 -584 9810
rect 584 9776 600 9810
rect -600 9729 600 9776
rect 658 9810 1858 9826
rect 658 9776 674 9810
rect 1842 9776 1858 9810
rect 658 9729 1858 9776
rect -1858 3303 -658 3329
rect -600 3303 600 3329
rect 658 3303 1858 3329
rect -1858 3245 -658 3261
rect -1858 3211 -1842 3245
rect -674 3211 -658 3245
rect -1858 3164 -658 3211
rect -600 3245 600 3261
rect -600 3211 -584 3245
rect 584 3211 600 3245
rect -600 3164 600 3211
rect 658 3245 1858 3261
rect 658 3211 674 3245
rect 1842 3211 1858 3245
rect 658 3164 1858 3211
rect -1858 -3262 -658 -3236
rect -600 -3262 600 -3236
rect 658 -3262 1858 -3236
rect -1858 -3320 -658 -3304
rect -1858 -3354 -1842 -3320
rect -674 -3354 -658 -3320
rect -1858 -3401 -658 -3354
rect -600 -3320 600 -3304
rect -600 -3354 -584 -3320
rect 584 -3354 600 -3320
rect -600 -3401 600 -3354
rect 658 -3320 1858 -3304
rect 658 -3354 674 -3320
rect 1842 -3354 1858 -3320
rect 658 -3401 1858 -3354
rect -1858 -9827 -658 -9801
rect -600 -9827 600 -9801
rect 658 -9827 1858 -9801
<< polycont >>
rect -1842 9776 -674 9810
rect -584 9776 584 9810
rect 674 9776 1842 9810
rect -1842 3211 -674 3245
rect -584 3211 584 3245
rect 674 3211 1842 3245
rect -1842 -3354 -674 -3320
rect -584 -3354 584 -3320
rect 674 -3354 1842 -3320
<< locali >>
rect -2038 9915 -1942 9949
rect 1942 9915 2038 9949
rect -2038 9853 -2004 9915
rect 2004 9853 2038 9915
rect -1858 9776 -1842 9810
rect -674 9776 -658 9810
rect -600 9776 -584 9810
rect 584 9776 600 9810
rect 658 9776 674 9810
rect 1842 9776 1858 9810
rect -1904 9717 -1870 9733
rect -1904 3325 -1870 3341
rect -646 9717 -612 9733
rect -646 3325 -612 3341
rect 612 9717 646 9733
rect 612 3325 646 3341
rect 1870 9717 1904 9733
rect 1870 3325 1904 3341
rect -1858 3211 -1842 3245
rect -674 3211 -658 3245
rect -600 3211 -584 3245
rect 584 3211 600 3245
rect 658 3211 674 3245
rect 1842 3211 1858 3245
rect -1904 3152 -1870 3168
rect -1904 -3240 -1870 -3224
rect -646 3152 -612 3168
rect -646 -3240 -612 -3224
rect 612 3152 646 3168
rect 612 -3240 646 -3224
rect 1870 3152 1904 3168
rect 1870 -3240 1904 -3224
rect -1858 -3354 -1842 -3320
rect -674 -3354 -658 -3320
rect -600 -3354 -584 -3320
rect 584 -3354 600 -3320
rect 658 -3354 674 -3320
rect 1842 -3354 1858 -3320
rect -1904 -3413 -1870 -3397
rect -1904 -9805 -1870 -9789
rect -646 -3413 -612 -3397
rect -646 -9805 -612 -9789
rect 612 -3413 646 -3397
rect 612 -9805 646 -9789
rect 1870 -3413 1904 -3397
rect 1870 -9805 1904 -9789
rect -2038 -9915 -2004 -9853
rect 2004 -9915 2038 -9853
rect -2038 -9949 -1942 -9915
rect 1942 -9949 2038 -9915
<< viali >>
rect -1842 9776 -674 9810
rect -584 9776 584 9810
rect 674 9776 1842 9810
rect -1904 3341 -1870 9717
rect -646 3341 -612 9717
rect 612 3341 646 9717
rect 1870 3341 1904 9717
rect -1842 3211 -674 3245
rect -584 3211 584 3245
rect 674 3211 1842 3245
rect -1904 -3224 -1870 3152
rect -646 -3224 -612 3152
rect 612 -3224 646 3152
rect 1870 -3224 1904 3152
rect -1842 -3354 -674 -3320
rect -584 -3354 584 -3320
rect 674 -3354 1842 -3320
rect -1904 -9789 -1870 -3413
rect -646 -9789 -612 -3413
rect 612 -9789 646 -3413
rect 1870 -9789 1904 -3413
<< metal1 >>
rect -1854 9810 -662 9816
rect -1854 9776 -1842 9810
rect -674 9776 -662 9810
rect -1854 9770 -662 9776
rect -596 9810 596 9816
rect -596 9776 -584 9810
rect 584 9776 596 9810
rect -596 9770 596 9776
rect 662 9810 1854 9816
rect 662 9776 674 9810
rect 1842 9776 1854 9810
rect 662 9770 1854 9776
rect -1910 9717 -1864 9729
rect -1910 3341 -1904 9717
rect -1870 3341 -1864 9717
rect -1910 3329 -1864 3341
rect -652 9717 -606 9729
rect -652 3341 -646 9717
rect -612 3341 -606 9717
rect -652 3329 -606 3341
rect 606 9717 652 9729
rect 606 3341 612 9717
rect 646 3341 652 9717
rect 606 3329 652 3341
rect 1864 9717 1910 9729
rect 1864 3341 1870 9717
rect 1904 3341 1910 9717
rect 1864 3329 1910 3341
rect -1854 3245 -662 3251
rect -1854 3211 -1842 3245
rect -674 3211 -662 3245
rect -1854 3205 -662 3211
rect -596 3245 596 3251
rect -596 3211 -584 3245
rect 584 3211 596 3245
rect -596 3205 596 3211
rect 662 3245 1854 3251
rect 662 3211 674 3245
rect 1842 3211 1854 3245
rect 662 3205 1854 3211
rect -1910 3152 -1864 3164
rect -1910 -3224 -1904 3152
rect -1870 -3224 -1864 3152
rect -1910 -3236 -1864 -3224
rect -652 3152 -606 3164
rect -652 -3224 -646 3152
rect -612 -3224 -606 3152
rect -652 -3236 -606 -3224
rect 606 3152 652 3164
rect 606 -3224 612 3152
rect 646 -3224 652 3152
rect 606 -3236 652 -3224
rect 1864 3152 1910 3164
rect 1864 -3224 1870 3152
rect 1904 -3224 1910 3152
rect 1864 -3236 1910 -3224
rect -1854 -3320 -662 -3314
rect -1854 -3354 -1842 -3320
rect -674 -3354 -662 -3320
rect -1854 -3360 -662 -3354
rect -596 -3320 596 -3314
rect -596 -3354 -584 -3320
rect 584 -3354 596 -3320
rect -596 -3360 596 -3354
rect 662 -3320 1854 -3314
rect 662 -3354 674 -3320
rect 1842 -3354 1854 -3320
rect 662 -3360 1854 -3354
rect -1910 -3413 -1864 -3401
rect -1910 -9789 -1904 -3413
rect -1870 -9789 -1864 -3413
rect -1910 -9801 -1864 -9789
rect -652 -3413 -606 -3401
rect -652 -9789 -646 -3413
rect -612 -9789 -606 -3413
rect -652 -9801 -606 -9789
rect 606 -3413 652 -3401
rect 606 -9789 612 -3413
rect 646 -9789 652 -3413
rect 606 -9801 652 -9789
rect 1864 -3413 1910 -3401
rect 1864 -9789 1870 -3413
rect 1904 -9789 1910 -3413
rect 1864 -9801 1910 -9789
<< properties >>
string FIXED_BBOX -2021 -9932 2021 9932
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 6.0 m 3 nf 3 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
