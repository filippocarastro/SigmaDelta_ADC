magic
tech sky130B
magscale 1 2
timestamp 1667069721
<< pwell >>
rect -828 -49239 828 49239
<< mvnmos >>
rect -600 39381 600 48981
rect -600 29563 600 39163
rect -600 19745 600 29345
rect -600 9927 600 19527
rect -600 109 600 9709
rect -600 -9709 600 -109
rect -600 -19527 600 -9927
rect -600 -29345 600 -19745
rect -600 -39163 600 -29563
rect -600 -48981 600 -39381
<< mvndiff >>
rect -658 48969 -600 48981
rect -658 39393 -646 48969
rect -612 39393 -600 48969
rect -658 39381 -600 39393
rect 600 48969 658 48981
rect 600 39393 612 48969
rect 646 39393 658 48969
rect 600 39381 658 39393
rect -658 39151 -600 39163
rect -658 29575 -646 39151
rect -612 29575 -600 39151
rect -658 29563 -600 29575
rect 600 39151 658 39163
rect 600 29575 612 39151
rect 646 29575 658 39151
rect 600 29563 658 29575
rect -658 29333 -600 29345
rect -658 19757 -646 29333
rect -612 19757 -600 29333
rect -658 19745 -600 19757
rect 600 29333 658 29345
rect 600 19757 612 29333
rect 646 19757 658 29333
rect 600 19745 658 19757
rect -658 19515 -600 19527
rect -658 9939 -646 19515
rect -612 9939 -600 19515
rect -658 9927 -600 9939
rect 600 19515 658 19527
rect 600 9939 612 19515
rect 646 9939 658 19515
rect 600 9927 658 9939
rect -658 9697 -600 9709
rect -658 121 -646 9697
rect -612 121 -600 9697
rect -658 109 -600 121
rect 600 9697 658 9709
rect 600 121 612 9697
rect 646 121 658 9697
rect 600 109 658 121
rect -658 -121 -600 -109
rect -658 -9697 -646 -121
rect -612 -9697 -600 -121
rect -658 -9709 -600 -9697
rect 600 -121 658 -109
rect 600 -9697 612 -121
rect 646 -9697 658 -121
rect 600 -9709 658 -9697
rect -658 -9939 -600 -9927
rect -658 -19515 -646 -9939
rect -612 -19515 -600 -9939
rect -658 -19527 -600 -19515
rect 600 -9939 658 -9927
rect 600 -19515 612 -9939
rect 646 -19515 658 -9939
rect 600 -19527 658 -19515
rect -658 -19757 -600 -19745
rect -658 -29333 -646 -19757
rect -612 -29333 -600 -19757
rect -658 -29345 -600 -29333
rect 600 -19757 658 -19745
rect 600 -29333 612 -19757
rect 646 -29333 658 -19757
rect 600 -29345 658 -29333
rect -658 -29575 -600 -29563
rect -658 -39151 -646 -29575
rect -612 -39151 -600 -29575
rect -658 -39163 -600 -39151
rect 600 -29575 658 -29563
rect 600 -39151 612 -29575
rect 646 -39151 658 -29575
rect 600 -39163 658 -39151
rect -658 -39393 -600 -39381
rect -658 -48969 -646 -39393
rect -612 -48969 -600 -39393
rect -658 -48981 -600 -48969
rect 600 -39393 658 -39381
rect 600 -48969 612 -39393
rect 646 -48969 658 -39393
rect 600 -48981 658 -48969
<< mvndiffc >>
rect -646 39393 -612 48969
rect 612 39393 646 48969
rect -646 29575 -612 39151
rect 612 29575 646 39151
rect -646 19757 -612 29333
rect 612 19757 646 29333
rect -646 9939 -612 19515
rect 612 9939 646 19515
rect -646 121 -612 9697
rect 612 121 646 9697
rect -646 -9697 -612 -121
rect 612 -9697 646 -121
rect -646 -19515 -612 -9939
rect 612 -19515 646 -9939
rect -646 -29333 -612 -19757
rect 612 -29333 646 -19757
rect -646 -39151 -612 -29575
rect 612 -39151 646 -29575
rect -646 -48969 -612 -39393
rect 612 -48969 646 -39393
<< mvpsubdiff >>
rect -792 49191 792 49203
rect -792 49157 -684 49191
rect 684 49157 792 49191
rect -792 49145 792 49157
rect -792 49095 -734 49145
rect -792 -49095 -780 49095
rect -746 -49095 -734 49095
rect 734 49095 792 49145
rect -792 -49145 -734 -49095
rect 734 -49095 746 49095
rect 780 -49095 792 49095
rect 734 -49145 792 -49095
rect -792 -49157 792 -49145
rect -792 -49191 -684 -49157
rect 684 -49191 792 -49157
rect -792 -49203 792 -49191
<< mvpsubdiffcont >>
rect -684 49157 684 49191
rect -780 -49095 -746 49095
rect 746 -49095 780 49095
rect -684 -49191 684 -49157
<< poly >>
rect -600 49053 600 49069
rect -600 49019 -584 49053
rect 584 49019 600 49053
rect -600 48981 600 49019
rect -600 39343 600 39381
rect -600 39309 -584 39343
rect 584 39309 600 39343
rect -600 39293 600 39309
rect -600 39235 600 39251
rect -600 39201 -584 39235
rect 584 39201 600 39235
rect -600 39163 600 39201
rect -600 29525 600 29563
rect -600 29491 -584 29525
rect 584 29491 600 29525
rect -600 29475 600 29491
rect -600 29417 600 29433
rect -600 29383 -584 29417
rect 584 29383 600 29417
rect -600 29345 600 29383
rect -600 19707 600 19745
rect -600 19673 -584 19707
rect 584 19673 600 19707
rect -600 19657 600 19673
rect -600 19599 600 19615
rect -600 19565 -584 19599
rect 584 19565 600 19599
rect -600 19527 600 19565
rect -600 9889 600 9927
rect -600 9855 -584 9889
rect 584 9855 600 9889
rect -600 9839 600 9855
rect -600 9781 600 9797
rect -600 9747 -584 9781
rect 584 9747 600 9781
rect -600 9709 600 9747
rect -600 71 600 109
rect -600 37 -584 71
rect 584 37 600 71
rect -600 21 600 37
rect -600 -37 600 -21
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -600 -109 600 -71
rect -600 -9747 600 -9709
rect -600 -9781 -584 -9747
rect 584 -9781 600 -9747
rect -600 -9797 600 -9781
rect -600 -9855 600 -9839
rect -600 -9889 -584 -9855
rect 584 -9889 600 -9855
rect -600 -9927 600 -9889
rect -600 -19565 600 -19527
rect -600 -19599 -584 -19565
rect 584 -19599 600 -19565
rect -600 -19615 600 -19599
rect -600 -19673 600 -19657
rect -600 -19707 -584 -19673
rect 584 -19707 600 -19673
rect -600 -19745 600 -19707
rect -600 -29383 600 -29345
rect -600 -29417 -584 -29383
rect 584 -29417 600 -29383
rect -600 -29433 600 -29417
rect -600 -29491 600 -29475
rect -600 -29525 -584 -29491
rect 584 -29525 600 -29491
rect -600 -29563 600 -29525
rect -600 -39201 600 -39163
rect -600 -39235 -584 -39201
rect 584 -39235 600 -39201
rect -600 -39251 600 -39235
rect -600 -39309 600 -39293
rect -600 -39343 -584 -39309
rect 584 -39343 600 -39309
rect -600 -39381 600 -39343
rect -600 -49019 600 -48981
rect -600 -49053 -584 -49019
rect 584 -49053 600 -49019
rect -600 -49069 600 -49053
<< polycont >>
rect -584 49019 584 49053
rect -584 39309 584 39343
rect -584 39201 584 39235
rect -584 29491 584 29525
rect -584 29383 584 29417
rect -584 19673 584 19707
rect -584 19565 584 19599
rect -584 9855 584 9889
rect -584 9747 584 9781
rect -584 37 584 71
rect -584 -71 584 -37
rect -584 -9781 584 -9747
rect -584 -9889 584 -9855
rect -584 -19599 584 -19565
rect -584 -19707 584 -19673
rect -584 -29417 584 -29383
rect -584 -29525 584 -29491
rect -584 -39235 584 -39201
rect -584 -39343 584 -39309
rect -584 -49053 584 -49019
<< locali >>
rect -780 49157 -684 49191
rect 684 49157 780 49191
rect -780 49095 -746 49157
rect 746 49095 780 49157
rect -600 49019 -584 49053
rect 584 49019 600 49053
rect -646 48969 -612 48985
rect -646 39377 -612 39393
rect 612 48969 646 48985
rect 612 39377 646 39393
rect -600 39309 -584 39343
rect 584 39309 600 39343
rect -600 39201 -584 39235
rect 584 39201 600 39235
rect -646 39151 -612 39167
rect -646 29559 -612 29575
rect 612 39151 646 39167
rect 612 29559 646 29575
rect -600 29491 -584 29525
rect 584 29491 600 29525
rect -600 29383 -584 29417
rect 584 29383 600 29417
rect -646 29333 -612 29349
rect -646 19741 -612 19757
rect 612 29333 646 29349
rect 612 19741 646 19757
rect -600 19673 -584 19707
rect 584 19673 600 19707
rect -600 19565 -584 19599
rect 584 19565 600 19599
rect -646 19515 -612 19531
rect -646 9923 -612 9939
rect 612 19515 646 19531
rect 612 9923 646 9939
rect -600 9855 -584 9889
rect 584 9855 600 9889
rect -600 9747 -584 9781
rect 584 9747 600 9781
rect -646 9697 -612 9713
rect -646 105 -612 121
rect 612 9697 646 9713
rect 612 105 646 121
rect -600 37 -584 71
rect 584 37 600 71
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -646 -121 -612 -105
rect -646 -9713 -612 -9697
rect 612 -121 646 -105
rect 612 -9713 646 -9697
rect -600 -9781 -584 -9747
rect 584 -9781 600 -9747
rect -600 -9889 -584 -9855
rect 584 -9889 600 -9855
rect -646 -9939 -612 -9923
rect -646 -19531 -612 -19515
rect 612 -9939 646 -9923
rect 612 -19531 646 -19515
rect -600 -19599 -584 -19565
rect 584 -19599 600 -19565
rect -600 -19707 -584 -19673
rect 584 -19707 600 -19673
rect -646 -19757 -612 -19741
rect -646 -29349 -612 -29333
rect 612 -19757 646 -19741
rect 612 -29349 646 -29333
rect -600 -29417 -584 -29383
rect 584 -29417 600 -29383
rect -600 -29525 -584 -29491
rect 584 -29525 600 -29491
rect -646 -29575 -612 -29559
rect -646 -39167 -612 -39151
rect 612 -29575 646 -29559
rect 612 -39167 646 -39151
rect -600 -39235 -584 -39201
rect 584 -39235 600 -39201
rect -600 -39343 -584 -39309
rect 584 -39343 600 -39309
rect -646 -39393 -612 -39377
rect -646 -48985 -612 -48969
rect 612 -39393 646 -39377
rect 612 -48985 646 -48969
rect -600 -49053 -584 -49019
rect 584 -49053 600 -49019
rect -780 -49157 -746 -49095
rect 746 -49157 780 -49095
rect -780 -49191 -684 -49157
rect 684 -49191 780 -49157
<< viali >>
rect -584 49019 584 49053
rect -646 39393 -612 48969
rect 612 39393 646 48969
rect -584 39309 584 39343
rect -584 39201 584 39235
rect -646 29575 -612 39151
rect 612 29575 646 39151
rect -584 29491 584 29525
rect -584 29383 584 29417
rect -646 19757 -612 29333
rect 612 19757 646 29333
rect -584 19673 584 19707
rect -584 19565 584 19599
rect -646 9939 -612 19515
rect 612 9939 646 19515
rect -584 9855 584 9889
rect -584 9747 584 9781
rect -646 121 -612 9697
rect 612 121 646 9697
rect -584 37 584 71
rect -584 -71 584 -37
rect -646 -9697 -612 -121
rect 612 -9697 646 -121
rect -584 -9781 584 -9747
rect -584 -9889 584 -9855
rect -646 -19515 -612 -9939
rect 612 -19515 646 -9939
rect -584 -19599 584 -19565
rect -584 -19707 584 -19673
rect -646 -29333 -612 -19757
rect 612 -29333 646 -19757
rect -584 -29417 584 -29383
rect -584 -29525 584 -29491
rect -646 -39151 -612 -29575
rect 612 -39151 646 -29575
rect -584 -39235 584 -39201
rect -584 -39343 584 -39309
rect -646 -48969 -612 -39393
rect 612 -48969 646 -39393
rect -584 -49053 584 -49019
<< metal1 >>
rect -596 49053 596 49059
rect -596 49019 -584 49053
rect 584 49019 596 49053
rect -596 49013 596 49019
rect -652 48969 -606 48981
rect -652 39393 -646 48969
rect -612 39393 -606 48969
rect -652 39381 -606 39393
rect 606 48969 652 48981
rect 606 39393 612 48969
rect 646 39393 652 48969
rect 606 39381 652 39393
rect -596 39343 596 39349
rect -596 39309 -584 39343
rect 584 39309 596 39343
rect -596 39303 596 39309
rect -596 39235 596 39241
rect -596 39201 -584 39235
rect 584 39201 596 39235
rect -596 39195 596 39201
rect -652 39151 -606 39163
rect -652 29575 -646 39151
rect -612 29575 -606 39151
rect -652 29563 -606 29575
rect 606 39151 652 39163
rect 606 29575 612 39151
rect 646 29575 652 39151
rect 606 29563 652 29575
rect -596 29525 596 29531
rect -596 29491 -584 29525
rect 584 29491 596 29525
rect -596 29485 596 29491
rect -596 29417 596 29423
rect -596 29383 -584 29417
rect 584 29383 596 29417
rect -596 29377 596 29383
rect -652 29333 -606 29345
rect -652 19757 -646 29333
rect -612 19757 -606 29333
rect -652 19745 -606 19757
rect 606 29333 652 29345
rect 606 19757 612 29333
rect 646 19757 652 29333
rect 606 19745 652 19757
rect -596 19707 596 19713
rect -596 19673 -584 19707
rect 584 19673 596 19707
rect -596 19667 596 19673
rect -596 19599 596 19605
rect -596 19565 -584 19599
rect 584 19565 596 19599
rect -596 19559 596 19565
rect -652 19515 -606 19527
rect -652 9939 -646 19515
rect -612 9939 -606 19515
rect -652 9927 -606 9939
rect 606 19515 652 19527
rect 606 9939 612 19515
rect 646 9939 652 19515
rect 606 9927 652 9939
rect -596 9889 596 9895
rect -596 9855 -584 9889
rect 584 9855 596 9889
rect -596 9849 596 9855
rect -596 9781 596 9787
rect -596 9747 -584 9781
rect 584 9747 596 9781
rect -596 9741 596 9747
rect -652 9697 -606 9709
rect -652 121 -646 9697
rect -612 121 -606 9697
rect -652 109 -606 121
rect 606 9697 652 9709
rect 606 121 612 9697
rect 646 121 652 9697
rect 606 109 652 121
rect -596 71 596 77
rect -596 37 -584 71
rect 584 37 596 71
rect -596 31 596 37
rect -596 -37 596 -31
rect -596 -71 -584 -37
rect 584 -71 596 -37
rect -596 -77 596 -71
rect -652 -121 -606 -109
rect -652 -9697 -646 -121
rect -612 -9697 -606 -121
rect -652 -9709 -606 -9697
rect 606 -121 652 -109
rect 606 -9697 612 -121
rect 646 -9697 652 -121
rect 606 -9709 652 -9697
rect -596 -9747 596 -9741
rect -596 -9781 -584 -9747
rect 584 -9781 596 -9747
rect -596 -9787 596 -9781
rect -596 -9855 596 -9849
rect -596 -9889 -584 -9855
rect 584 -9889 596 -9855
rect -596 -9895 596 -9889
rect -652 -9939 -606 -9927
rect -652 -19515 -646 -9939
rect -612 -19515 -606 -9939
rect -652 -19527 -606 -19515
rect 606 -9939 652 -9927
rect 606 -19515 612 -9939
rect 646 -19515 652 -9939
rect 606 -19527 652 -19515
rect -596 -19565 596 -19559
rect -596 -19599 -584 -19565
rect 584 -19599 596 -19565
rect -596 -19605 596 -19599
rect -596 -19673 596 -19667
rect -596 -19707 -584 -19673
rect 584 -19707 596 -19673
rect -596 -19713 596 -19707
rect -652 -19757 -606 -19745
rect -652 -29333 -646 -19757
rect -612 -29333 -606 -19757
rect -652 -29345 -606 -29333
rect 606 -19757 652 -19745
rect 606 -29333 612 -19757
rect 646 -29333 652 -19757
rect 606 -29345 652 -29333
rect -596 -29383 596 -29377
rect -596 -29417 -584 -29383
rect 584 -29417 596 -29383
rect -596 -29423 596 -29417
rect -596 -29491 596 -29485
rect -596 -29525 -584 -29491
rect 584 -29525 596 -29491
rect -596 -29531 596 -29525
rect -652 -29575 -606 -29563
rect -652 -39151 -646 -29575
rect -612 -39151 -606 -29575
rect -652 -39163 -606 -39151
rect 606 -29575 652 -29563
rect 606 -39151 612 -29575
rect 646 -39151 652 -29575
rect 606 -39163 652 -39151
rect -596 -39201 596 -39195
rect -596 -39235 -584 -39201
rect 584 -39235 596 -39201
rect -596 -39241 596 -39235
rect -596 -39309 596 -39303
rect -596 -39343 -584 -39309
rect 584 -39343 596 -39309
rect -596 -39349 596 -39343
rect -652 -39393 -606 -39381
rect -652 -48969 -646 -39393
rect -612 -48969 -606 -39393
rect -652 -48981 -606 -48969
rect 606 -39393 652 -39381
rect 606 -48969 612 -39393
rect 646 -48969 652 -39393
rect 606 -48981 652 -48969
rect -596 -49019 596 -49013
rect -596 -49053 -584 -49019
rect 584 -49053 596 -49019
rect -596 -49059 596 -49053
<< properties >>
string FIXED_BBOX -763 -49174 763 49174
string gencell sky130_fd_pr__nfet_g5v0d10v5
string library sky130
string parameters w 48.0 l 6.0 m 10 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
