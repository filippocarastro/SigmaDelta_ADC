magic
tech sky130B
magscale 1 2
timestamp 1667656102
<< metal1 >>
rect 38942 36638 39422 36642
rect 11988 35104 44904 36638
rect 11988 35102 42004 35104
rect 42778 35102 44904 35104
rect 14754 30634 15404 35102
rect 16160 30742 16768 34724
rect 16160 30534 16342 30742
rect 16578 30534 16768 30742
rect 17416 30642 18066 35102
rect 18676 30742 19284 34742
rect 16160 30452 16768 30534
rect 18676 30534 18848 30742
rect 19084 30534 19284 30742
rect 19868 30652 20518 35102
rect 21174 30760 21782 34760
rect 18676 30470 19284 30534
rect 21174 30552 21346 30760
rect 21582 30552 21782 30760
rect 22374 30652 23024 35102
rect 23708 30742 24316 34770
rect 21174 30488 21782 30552
rect 23708 30534 23880 30742
rect 24116 30534 24316 30742
rect 24882 30652 25532 35102
rect 26214 30742 26822 34742
rect 23708 30498 24316 30534
rect 26214 30534 26396 30742
rect 26632 30534 26822 30742
rect 27406 30642 28056 35102
rect 28722 30732 29330 34760
rect 26214 30470 26822 30534
rect 28722 30524 28894 30732
rect 29130 30524 29330 30732
rect 29912 30652 30562 35102
rect 31228 30768 31836 34788
rect 28722 30488 29330 30524
rect 31228 30560 31418 30768
rect 31654 30560 31836 30768
rect 32446 30652 33096 35102
rect 33744 30742 34352 34770
rect 31228 30516 31836 30560
rect 33744 30534 33934 30742
rect 34170 30534 34352 30742
rect 35100 30655 35750 35102
rect 36402 30676 36882 35102
rect 37688 31140 38170 34784
rect 37688 30914 37786 31140
rect 38066 30914 38170 31140
rect 37688 30768 38170 30914
rect 38942 30706 39422 35102
rect 40190 31104 40672 34816
rect 40190 30878 40274 31104
rect 40554 30878 40672 31104
rect 40190 30800 40672 30878
rect 41524 30702 42004 35102
rect 42378 34378 42752 34680
rect 33744 30498 34352 30534
rect 14835 30290 37650 30291
rect 42378 30290 42680 34378
rect 43912 30614 44884 35102
rect 14835 30287 43690 30290
rect 14835 30248 43857 30287
rect 14835 29801 43858 30248
rect 14835 29499 45329 29801
rect 14835 29406 43858 29499
rect 14835 29404 43690 29406
rect 13848 28028 14048 28228
rect 26604 28092 34477 28498
rect 35227 28214 35813 28343
rect 35227 28002 35394 28214
rect 35590 28002 35813 28214
rect 36758 28190 45408 28602
rect 14777 25544 24229 25846
rect 14976 25388 15610 25438
rect 14976 25188 15190 25388
rect 15390 25188 15610 25388
rect 13316 16036 14520 24924
rect 14976 16984 15610 25188
rect 17548 25400 18182 25426
rect 17548 25200 17808 25400
rect 18008 25200 18182 25400
rect 16176 16036 16924 24860
rect 17548 16972 18182 25200
rect 20736 25226 21472 25234
rect 18716 16036 19464 24872
rect 19882 24490 20736 24748
rect 19882 24294 21472 24490
rect 23927 24360 24229 25544
rect 23926 24354 24230 24360
rect 19882 23896 21428 24294
rect 21826 23896 21832 24294
rect 23926 24044 24230 24050
rect 19882 16632 21472 23896
rect 27514 21634 28100 27878
rect 27514 21390 27644 21634
rect 27886 21390 28100 21634
rect 28915 22245 29581 27827
rect 30122 22568 30642 27850
rect 30122 22394 30324 22568
rect 30524 22394 30642 22568
rect 30122 22312 30642 22394
rect 31375 22245 32041 27791
rect 32682 22596 33202 27896
rect 32682 22422 32846 22596
rect 33046 22422 33202 22596
rect 32682 22358 33202 22422
rect 34092 27847 34678 27848
rect 35227 27847 35813 28002
rect 37368 28030 37860 28082
rect 34092 27261 35813 27847
rect 34092 22245 34678 27261
rect 28915 21579 34678 22245
rect 36006 22496 36482 27922
rect 37368 27830 37524 28030
rect 37724 27830 37860 28030
rect 39882 28030 40374 28090
rect 37368 22594 37860 27830
rect 38626 22496 39102 27902
rect 39882 27830 40046 28030
rect 40246 27830 40374 28030
rect 42402 28038 42894 28120
rect 39882 22602 40374 27830
rect 41144 22496 41620 27902
rect 42402 27838 42542 28038
rect 42742 27838 42894 28038
rect 42402 22632 42894 27838
rect 43766 22496 44222 27916
rect 36006 22020 44222 22496
rect 27514 21206 28100 21390
rect 27514 20844 43715 21206
rect 27514 16551 28100 20844
rect 28908 16036 29454 20420
rect 41680 16593 42648 20404
rect 43766 16860 44222 22020
rect 41680 16036 42661 16593
rect 43766 16404 44914 16860
rect 45370 16404 45376 16860
rect 43766 16198 44222 16404
rect 11752 16014 43830 16036
rect 11752 13988 45222 16014
<< via1 >>
rect 16342 30534 16578 30742
rect 18848 30534 19084 30742
rect 21346 30552 21582 30760
rect 23880 30534 24116 30742
rect 26396 30534 26632 30742
rect 28894 30524 29130 30732
rect 31418 30560 31654 30768
rect 33934 30534 34170 30742
rect 37786 30914 38066 31140
rect 40274 30878 40554 31104
rect 35394 28002 35590 28214
rect 15190 25188 15390 25388
rect 17808 25200 18008 25400
rect 20736 24490 21472 25226
rect 21428 23896 21826 24294
rect 23926 24050 24230 24354
rect 27644 21390 27886 21634
rect 30324 22394 30524 22568
rect 32846 22422 33046 22596
rect 37524 27830 37724 28030
rect 40046 27830 40246 28030
rect 42542 27838 42742 28038
rect 44914 16404 45370 16860
<< metal2 >>
rect 35918 31140 40800 31249
rect 35918 30914 37786 31140
rect 38066 31104 40800 31140
rect 38066 30914 40274 31104
rect 13560 30768 34904 30910
rect 13560 30760 31418 30768
rect 13560 30742 21346 30760
rect 13560 30534 16342 30742
rect 16578 30534 18848 30742
rect 19084 30552 21346 30742
rect 21582 30742 31418 30760
rect 21582 30552 23880 30742
rect 19084 30534 23880 30552
rect 24116 30534 26396 30742
rect 26632 30732 31418 30742
rect 26632 30534 28894 30732
rect 13560 30524 28894 30534
rect 29130 30560 31418 30732
rect 31654 30742 34904 30768
rect 31654 30560 33934 30742
rect 29130 30534 33934 30560
rect 34170 30534 34904 30742
rect 29130 30524 34904 30534
rect 13560 30173 34904 30524
rect 35918 30878 40274 30914
rect 40554 30878 40800 31104
rect 35918 30716 40800 30878
rect 13560 28435 14297 30173
rect 35918 29443 36451 30716
rect 35286 28910 36451 29443
rect 13560 27698 21473 28435
rect 35286 28303 35798 28910
rect 35286 28214 43508 28303
rect 35286 28002 35394 28214
rect 35590 28038 43508 28214
rect 35590 28030 42542 28038
rect 35590 28002 37524 28030
rect 35286 27830 37524 28002
rect 37724 27830 40046 28030
rect 40246 27838 42542 28030
rect 42742 27838 43508 28038
rect 40246 27830 43508 27838
rect 35286 27770 43508 27830
rect 20736 25438 21472 27698
rect 14794 25400 21472 25438
rect 14794 25388 17808 25400
rect 14794 25188 15190 25388
rect 15390 25200 17808 25388
rect 18008 25226 21472 25400
rect 18008 25200 20736 25226
rect 15390 25188 20736 25200
rect 14794 25006 20736 25188
rect 20730 24490 20736 25006
rect 21472 24490 21478 25226
rect 21428 24294 21826 24300
rect 21826 23896 22053 24294
rect 22451 23896 22460 24294
rect 23920 24050 23926 24354
rect 24230 24050 24236 24354
rect 21428 23890 21826 23896
rect 23926 20950 24230 24050
rect 28071 22596 33741 22623
rect 28071 22568 32846 22596
rect 28071 22394 30324 22568
rect 30524 22422 32846 22568
rect 33046 22422 33741 22596
rect 30524 22394 33741 22422
rect 28071 22037 33741 22394
rect 28071 21876 28657 22037
rect 28176 21726 28657 21876
rect 27512 21634 28657 21726
rect 27512 21390 27644 21634
rect 27886 21390 28657 21634
rect 27512 21245 28657 21390
rect 23742 20550 24230 20950
rect 23742 16860 24198 20550
rect 44914 16860 45370 16866
rect 23742 16404 44914 16860
rect 44914 16398 45370 16404
<< via2 >>
rect 22053 23896 22451 24294
<< metal3 >>
rect 22048 24294 22456 24299
rect 22048 23896 22053 24294
rect 22451 23896 23310 24294
rect 22048 23891 22456 23896
rect 22643 23666 23310 23896
rect 22642 22692 23310 23666
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1667223724
transform 1 0 24090 0 1 20400
box -3150 -3100 3149 3100
use sky130_fd_pr__nfet_g5v0d10v5_U4FG9E  XM1
timestamp 1667224822
transform 1 0 43184 0 1 18477
box -828 -2627 828 2627
use sky130_fd_pr__pfet_g5v0d10v5_VS8EJU  XM2
timestamp 1667224016
transform 1 0 31046 0 -1 25238
box -3374 -3462 3374 3462
use sky130_fd_pr__nfet_01v8_45ERJ4  XM3
timestamp 1667324858
transform 1 0 28674 0 1 18483
box -796 -2579 796 2579
use sky130_fd_pr__pfet_g5v0d10v5_VS8V9Y  XM4
timestamp 1667223724
transform 1 0 40119 0 1 25266
box -4003 -3462 4003 3462
use sky130_fd_pr__pfet_g5v0d10v5_VSGFLU  XM5
timestamp 1667223724
transform -1 0 39185 0 -1 32696
box -2745 -2662 2745 2662
use sky130_fd_pr__pfet_g5v0d10v5_YHBQGB  XM6
timestamp 1667223724
transform 1 0 25251 0 1 32660
box -10293 -2662 10293 2662
use sky130_fd_pr__nfet_g5v0d10v5_8VPWNZ  XM7
timestamp 1667325532
transform 1 0 17202 0 1 20921
box -3344 -5027 3344 5027
use sky130_fd_pr__pfet_g5v0d10v5_VSGNQY  XM8
timestamp 1667223724
transform 1 0 43332 0 1 32694
box -858 -2662 858 2662
<< labels >>
flabel metal1 12642 35948 12842 36148 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 45106 29566 45306 29766 0 FreeSans 256 0 0 0 Ibias
port 4 nsew
flabel metal1 45192 28196 45392 28396 0 FreeSans 256 0 0 0 Vinp
port 1 nsew
flabel metal1 26604 28092 26804 28292 0 FreeSans 256 0 0 0 Vinn
port 0 nsew
flabel metal1 44802 14338 45002 14538 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 13848 28028 14048 28228 0 FreeSans 256 0 0 0 Vout
port 5 nsew
<< end >>
