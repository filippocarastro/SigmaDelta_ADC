magic
tech sky130B
magscale 1 2
timestamp 1667120857
<< nwell >>
rect -2745 -6744 2745 6744
<< mvpmos >>
rect -2487 47 -1287 6447
rect -1229 47 -29 6447
rect 29 47 1229 6447
rect 1287 47 2487 6447
rect -2487 -6518 -1287 -118
rect -1229 -6518 -29 -118
rect 29 -6518 1229 -118
rect 1287 -6518 2487 -118
<< mvpdiff >>
rect -2545 6435 -2487 6447
rect -2545 59 -2533 6435
rect -2499 59 -2487 6435
rect -2545 47 -2487 59
rect -1287 6435 -1229 6447
rect -1287 59 -1275 6435
rect -1241 59 -1229 6435
rect -1287 47 -1229 59
rect -29 6435 29 6447
rect -29 59 -17 6435
rect 17 59 29 6435
rect -29 47 29 59
rect 1229 6435 1287 6447
rect 1229 59 1241 6435
rect 1275 59 1287 6435
rect 1229 47 1287 59
rect 2487 6435 2545 6447
rect 2487 59 2499 6435
rect 2533 59 2545 6435
rect 2487 47 2545 59
rect -2545 -130 -2487 -118
rect -2545 -6506 -2533 -130
rect -2499 -6506 -2487 -130
rect -2545 -6518 -2487 -6506
rect -1287 -130 -1229 -118
rect -1287 -6506 -1275 -130
rect -1241 -6506 -1229 -130
rect -1287 -6518 -1229 -6506
rect -29 -130 29 -118
rect -29 -6506 -17 -130
rect 17 -6506 29 -130
rect -29 -6518 29 -6506
rect 1229 -130 1287 -118
rect 1229 -6506 1241 -130
rect 1275 -6506 1287 -130
rect 1229 -6518 1287 -6506
rect 2487 -130 2545 -118
rect 2487 -6506 2499 -130
rect 2533 -6506 2545 -130
rect 2487 -6518 2545 -6506
<< mvpdiffc >>
rect -2533 59 -2499 6435
rect -1275 59 -1241 6435
rect -17 59 17 6435
rect 1241 59 1275 6435
rect 2499 59 2533 6435
rect -2533 -6506 -2499 -130
rect -1275 -6506 -1241 -130
rect -17 -6506 17 -130
rect 1241 -6506 1275 -130
rect 2499 -6506 2533 -130
<< mvnsubdiff >>
rect -2679 6666 2679 6678
rect -2679 6632 -2571 6666
rect 2571 6632 2679 6666
rect -2679 6620 2679 6632
rect -2679 6570 -2621 6620
rect -2679 -6570 -2667 6570
rect -2633 -6570 -2621 6570
rect 2621 6570 2679 6620
rect -2679 -6620 -2621 -6570
rect 2621 -6570 2633 6570
rect 2667 -6570 2679 6570
rect 2621 -6620 2679 -6570
rect -2679 -6632 2679 -6620
rect -2679 -6666 -2571 -6632
rect 2571 -6666 2679 -6632
rect -2679 -6678 2679 -6666
<< mvnsubdiffcont >>
rect -2571 6632 2571 6666
rect -2667 -6570 -2633 6570
rect 2633 -6570 2667 6570
rect -2571 -6666 2571 -6632
<< poly >>
rect -2487 6528 -1287 6544
rect -2487 6494 -2471 6528
rect -1303 6494 -1287 6528
rect -2487 6447 -1287 6494
rect -1229 6528 -29 6544
rect -1229 6494 -1213 6528
rect -45 6494 -29 6528
rect -1229 6447 -29 6494
rect 29 6528 1229 6544
rect 29 6494 45 6528
rect 1213 6494 1229 6528
rect 29 6447 1229 6494
rect 1287 6528 2487 6544
rect 1287 6494 1303 6528
rect 2471 6494 2487 6528
rect 1287 6447 2487 6494
rect -2487 21 -1287 47
rect -1229 21 -29 47
rect 29 21 1229 47
rect 1287 21 2487 47
rect -2487 -37 -1287 -21
rect -2487 -71 -2471 -37
rect -1303 -71 -1287 -37
rect -2487 -118 -1287 -71
rect -1229 -37 -29 -21
rect -1229 -71 -1213 -37
rect -45 -71 -29 -37
rect -1229 -118 -29 -71
rect 29 -37 1229 -21
rect 29 -71 45 -37
rect 1213 -71 1229 -37
rect 29 -118 1229 -71
rect 1287 -37 2487 -21
rect 1287 -71 1303 -37
rect 2471 -71 2487 -37
rect 1287 -118 2487 -71
rect -2487 -6544 -1287 -6518
rect -1229 -6544 -29 -6518
rect 29 -6544 1229 -6518
rect 1287 -6544 2487 -6518
<< polycont >>
rect -2471 6494 -1303 6528
rect -1213 6494 -45 6528
rect 45 6494 1213 6528
rect 1303 6494 2471 6528
rect -2471 -71 -1303 -37
rect -1213 -71 -45 -37
rect 45 -71 1213 -37
rect 1303 -71 2471 -37
<< locali >>
rect -2667 6632 -2571 6666
rect 2571 6632 2667 6666
rect -2667 6570 -2633 6632
rect 2633 6570 2667 6632
rect -2487 6494 -2471 6528
rect -1303 6494 -1287 6528
rect -1229 6494 -1213 6528
rect -45 6494 -29 6528
rect 29 6494 45 6528
rect 1213 6494 1229 6528
rect 1287 6494 1303 6528
rect 2471 6494 2487 6528
rect -2533 6435 -2499 6451
rect -2533 43 -2499 59
rect -1275 6435 -1241 6451
rect -1275 43 -1241 59
rect -17 6435 17 6451
rect -17 43 17 59
rect 1241 6435 1275 6451
rect 1241 43 1275 59
rect 2499 6435 2533 6451
rect 2499 43 2533 59
rect -2487 -71 -2471 -37
rect -1303 -71 -1287 -37
rect -1229 -71 -1213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1213 -71 1229 -37
rect 1287 -71 1303 -37
rect 2471 -71 2487 -37
rect -2533 -130 -2499 -114
rect -2533 -6522 -2499 -6506
rect -1275 -130 -1241 -114
rect -1275 -6522 -1241 -6506
rect -17 -130 17 -114
rect -17 -6522 17 -6506
rect 1241 -130 1275 -114
rect 1241 -6522 1275 -6506
rect 2499 -130 2533 -114
rect 2499 -6522 2533 -6506
rect -2667 -6632 -2633 -6570
rect 2633 -6632 2667 -6570
rect -2667 -6666 -2571 -6632
rect 2571 -6666 2667 -6632
<< viali >>
rect -2471 6494 -1303 6528
rect -1213 6494 -45 6528
rect 45 6494 1213 6528
rect 1303 6494 2471 6528
rect -2533 59 -2499 6435
rect -1275 59 -1241 6435
rect -17 59 17 6435
rect 1241 59 1275 6435
rect 2499 59 2533 6435
rect -2471 -71 -1303 -37
rect -1213 -71 -45 -37
rect 45 -71 1213 -37
rect 1303 -71 2471 -37
rect -2533 -6506 -2499 -130
rect -1275 -6506 -1241 -130
rect -17 -6506 17 -130
rect 1241 -6506 1275 -130
rect 2499 -6506 2533 -130
<< metal1 >>
rect -2483 6528 -1291 6534
rect -2483 6494 -2471 6528
rect -1303 6494 -1291 6528
rect -2483 6488 -1291 6494
rect -1225 6528 -33 6534
rect -1225 6494 -1213 6528
rect -45 6494 -33 6528
rect -1225 6488 -33 6494
rect 33 6528 1225 6534
rect 33 6494 45 6528
rect 1213 6494 1225 6528
rect 33 6488 1225 6494
rect 1291 6528 2483 6534
rect 1291 6494 1303 6528
rect 2471 6494 2483 6528
rect 1291 6488 2483 6494
rect -2539 6435 -2493 6447
rect -2539 59 -2533 6435
rect -2499 59 -2493 6435
rect -2539 47 -2493 59
rect -1281 6435 -1235 6447
rect -1281 59 -1275 6435
rect -1241 59 -1235 6435
rect -1281 47 -1235 59
rect -23 6435 23 6447
rect -23 59 -17 6435
rect 17 59 23 6435
rect -23 47 23 59
rect 1235 6435 1281 6447
rect 1235 59 1241 6435
rect 1275 59 1281 6435
rect 1235 47 1281 59
rect 2493 6435 2539 6447
rect 2493 59 2499 6435
rect 2533 59 2539 6435
rect 2493 47 2539 59
rect -2483 -37 -1291 -31
rect -2483 -71 -2471 -37
rect -1303 -71 -1291 -37
rect -2483 -77 -1291 -71
rect -1225 -37 -33 -31
rect -1225 -71 -1213 -37
rect -45 -71 -33 -37
rect -1225 -77 -33 -71
rect 33 -37 1225 -31
rect 33 -71 45 -37
rect 1213 -71 1225 -37
rect 33 -77 1225 -71
rect 1291 -37 2483 -31
rect 1291 -71 1303 -37
rect 2471 -71 2483 -37
rect 1291 -77 2483 -71
rect -2539 -130 -2493 -118
rect -2539 -6506 -2533 -130
rect -2499 -6506 -2493 -130
rect -2539 -6518 -2493 -6506
rect -1281 -130 -1235 -118
rect -1281 -6506 -1275 -130
rect -1241 -6506 -1235 -130
rect -1281 -6518 -1235 -6506
rect -23 -130 23 -118
rect -23 -6506 -17 -130
rect 17 -6506 23 -130
rect -23 -6518 23 -6506
rect 1235 -130 1281 -118
rect 1235 -6506 1241 -130
rect 1275 -6506 1281 -130
rect 1235 -6518 1281 -6506
rect 2493 -130 2539 -118
rect 2493 -6506 2499 -130
rect 2533 -6506 2539 -130
rect 2493 -6518 2539 -6506
<< properties >>
string FIXED_BBOX -2650 -6649 2650 6649
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 6.0 m 2 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
