magic
tech sky130B
magscale 1 2
timestamp 1667211484
<< metal1 >>
rect 11988 35104 44904 36638
rect 11988 35102 41536 35104
rect 42778 35102 44904 35104
rect 43912 30614 44884 35102
rect 42806 30248 43856 30284
rect 42806 29764 43858 30248
rect 16562 25252 16762 25452
rect 12828 6758 13028 6958
rect 14266 6710 14466 6910
rect 15146 6706 15346 6906
rect 16380 6638 16580 6838
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1667069721
transform 1 0 15164 0 1 14122
box -3150 -3100 3149 3100
use sky130_fd_pr__nfet_g5v0d10v5_S447FE  XM1
timestamp 1667069824
transform 1 0 26542 0 1 13409
box -828 -2627 828 2627
use sky130_fd_pr__pfet_g5v0d10v5_AGKGBY  XM2
timestamp 1667120857
transform 1 0 36618 0 -1 25490
box -3374 -3462 3374 3462
use sky130_fd_pr__nfet_01v8_B39JSP  XM3
timestamp 1667121247
transform 1 0 20618 0 1 13601
box -796 -2579 796 2579
use sky130_fd_pr__pfet_g5v0d10v5_AGFYAY  XM4
timestamp 1667069824
transform 1 0 23335 0 1 25352
box -4003 -3462 4003 3462
use sky130_fd_pr__pfet_g5v0d10v5_NGD7BL  XM5
timestamp 1667120857
transform -1 0 15191 0 -1 32732
box -2745 -2662 2745 2662
use sky130_fd_pr__pfet_g5v0d10v5_PEV8FT  XM6
timestamp 1667069824
transform 1 0 29619 0 1 32754
box -10293 -2662 10293 2662
use sky130_fd_pr__nfet_g5v0d10v5_59B6FY  XM7
timestamp 1667069824
transform 1 0 36772 0 1 15917
box -3344 -5027 3344 5027
use sky130_fd_pr__pfet_g5v0d10v5_VSGNQY  XM8
timestamp 1667211103
transform 1 0 43332 0 1 32694
box -858 -2662 858 2662
<< labels >>
flabel metal1 16562 25252 16762 25452 0 FreeSans 256 0 0 0 Vinn
port 0 nsew
flabel metal1 12642 35948 12842 36148 0 FreeSans 256 0 0 0 VDD
port 3 nsew
flabel metal1 12828 6758 13028 6958 0 FreeSans 256 0 0 0 Vinp
port 1 nsew
flabel metal1 14266 6710 14466 6910 0 FreeSans 256 0 0 0 GND
port 2 nsew
flabel metal1 15146 6706 15346 6906 0 FreeSans 256 0 0 0 Vout
port 5 nsew
flabel metal1 16380 6638 16580 6838 0 FreeSans 256 0 0 0 Ibias
port 4 nsew
<< end >>
