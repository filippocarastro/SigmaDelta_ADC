magic
tech sky130B
magscale 1 2
timestamp 1667069721
<< nwell >>
rect -2745 -10251 2745 10251
<< mvpmos >>
rect -2487 5154 -1287 9954
rect -1229 5154 -29 9954
rect 29 5154 1229 9954
rect 1287 5154 2487 9954
rect -2487 118 -1287 4918
rect -1229 118 -29 4918
rect 29 118 1229 4918
rect 1287 118 2487 4918
rect -2487 -4918 -1287 -118
rect -1229 -4918 -29 -118
rect 29 -4918 1229 -118
rect 1287 -4918 2487 -118
rect -2487 -9954 -1287 -5154
rect -1229 -9954 -29 -5154
rect 29 -9954 1229 -5154
rect 1287 -9954 2487 -5154
<< mvpdiff >>
rect -2545 9942 -2487 9954
rect -2545 5166 -2533 9942
rect -2499 5166 -2487 9942
rect -2545 5154 -2487 5166
rect -1287 9942 -1229 9954
rect -1287 5166 -1275 9942
rect -1241 5166 -1229 9942
rect -1287 5154 -1229 5166
rect -29 9942 29 9954
rect -29 5166 -17 9942
rect 17 5166 29 9942
rect -29 5154 29 5166
rect 1229 9942 1287 9954
rect 1229 5166 1241 9942
rect 1275 5166 1287 9942
rect 1229 5154 1287 5166
rect 2487 9942 2545 9954
rect 2487 5166 2499 9942
rect 2533 5166 2545 9942
rect 2487 5154 2545 5166
rect -2545 4906 -2487 4918
rect -2545 130 -2533 4906
rect -2499 130 -2487 4906
rect -2545 118 -2487 130
rect -1287 4906 -1229 4918
rect -1287 130 -1275 4906
rect -1241 130 -1229 4906
rect -1287 118 -1229 130
rect -29 4906 29 4918
rect -29 130 -17 4906
rect 17 130 29 4906
rect -29 118 29 130
rect 1229 4906 1287 4918
rect 1229 130 1241 4906
rect 1275 130 1287 4906
rect 1229 118 1287 130
rect 2487 4906 2545 4918
rect 2487 130 2499 4906
rect 2533 130 2545 4906
rect 2487 118 2545 130
rect -2545 -130 -2487 -118
rect -2545 -4906 -2533 -130
rect -2499 -4906 -2487 -130
rect -2545 -4918 -2487 -4906
rect -1287 -130 -1229 -118
rect -1287 -4906 -1275 -130
rect -1241 -4906 -1229 -130
rect -1287 -4918 -1229 -4906
rect -29 -130 29 -118
rect -29 -4906 -17 -130
rect 17 -4906 29 -130
rect -29 -4918 29 -4906
rect 1229 -130 1287 -118
rect 1229 -4906 1241 -130
rect 1275 -4906 1287 -130
rect 1229 -4918 1287 -4906
rect 2487 -130 2545 -118
rect 2487 -4906 2499 -130
rect 2533 -4906 2545 -130
rect 2487 -4918 2545 -4906
rect -2545 -5166 -2487 -5154
rect -2545 -9942 -2533 -5166
rect -2499 -9942 -2487 -5166
rect -2545 -9954 -2487 -9942
rect -1287 -5166 -1229 -5154
rect -1287 -9942 -1275 -5166
rect -1241 -9942 -1229 -5166
rect -1287 -9954 -1229 -9942
rect -29 -5166 29 -5154
rect -29 -9942 -17 -5166
rect 17 -9942 29 -5166
rect -29 -9954 29 -9942
rect 1229 -5166 1287 -5154
rect 1229 -9942 1241 -5166
rect 1275 -9942 1287 -5166
rect 1229 -9954 1287 -9942
rect 2487 -5166 2545 -5154
rect 2487 -9942 2499 -5166
rect 2533 -9942 2545 -5166
rect 2487 -9954 2545 -9942
<< mvpdiffc >>
rect -2533 5166 -2499 9942
rect -1275 5166 -1241 9942
rect -17 5166 17 9942
rect 1241 5166 1275 9942
rect 2499 5166 2533 9942
rect -2533 130 -2499 4906
rect -1275 130 -1241 4906
rect -17 130 17 4906
rect 1241 130 1275 4906
rect 2499 130 2533 4906
rect -2533 -4906 -2499 -130
rect -1275 -4906 -1241 -130
rect -17 -4906 17 -130
rect 1241 -4906 1275 -130
rect 2499 -4906 2533 -130
rect -2533 -9942 -2499 -5166
rect -1275 -9942 -1241 -5166
rect -17 -9942 17 -5166
rect 1241 -9942 1275 -5166
rect 2499 -9942 2533 -5166
<< mvnsubdiff >>
rect -2679 10173 2679 10185
rect -2679 10139 -2571 10173
rect 2571 10139 2679 10173
rect -2679 10127 2679 10139
rect -2679 10077 -2621 10127
rect -2679 -10077 -2667 10077
rect -2633 -10077 -2621 10077
rect 2621 10077 2679 10127
rect -2679 -10127 -2621 -10077
rect 2621 -10077 2633 10077
rect 2667 -10077 2679 10077
rect 2621 -10127 2679 -10077
rect -2679 -10139 2679 -10127
rect -2679 -10173 -2571 -10139
rect 2571 -10173 2679 -10139
rect -2679 -10185 2679 -10173
<< mvnsubdiffcont >>
rect -2571 10139 2571 10173
rect -2667 -10077 -2633 10077
rect 2633 -10077 2667 10077
rect -2571 -10173 2571 -10139
<< poly >>
rect -2487 10035 -1287 10051
rect -2487 10001 -2471 10035
rect -1303 10001 -1287 10035
rect -2487 9954 -1287 10001
rect -1229 10035 -29 10051
rect -1229 10001 -1213 10035
rect -45 10001 -29 10035
rect -1229 9954 -29 10001
rect 29 10035 1229 10051
rect 29 10001 45 10035
rect 1213 10001 1229 10035
rect 29 9954 1229 10001
rect 1287 10035 2487 10051
rect 1287 10001 1303 10035
rect 2471 10001 2487 10035
rect 1287 9954 2487 10001
rect -2487 5107 -1287 5154
rect -2487 5073 -2471 5107
rect -1303 5073 -1287 5107
rect -2487 5057 -1287 5073
rect -1229 5107 -29 5154
rect -1229 5073 -1213 5107
rect -45 5073 -29 5107
rect -1229 5057 -29 5073
rect 29 5107 1229 5154
rect 29 5073 45 5107
rect 1213 5073 1229 5107
rect 29 5057 1229 5073
rect 1287 5107 2487 5154
rect 1287 5073 1303 5107
rect 2471 5073 2487 5107
rect 1287 5057 2487 5073
rect -2487 4999 -1287 5015
rect -2487 4965 -2471 4999
rect -1303 4965 -1287 4999
rect -2487 4918 -1287 4965
rect -1229 4999 -29 5015
rect -1229 4965 -1213 4999
rect -45 4965 -29 4999
rect -1229 4918 -29 4965
rect 29 4999 1229 5015
rect 29 4965 45 4999
rect 1213 4965 1229 4999
rect 29 4918 1229 4965
rect 1287 4999 2487 5015
rect 1287 4965 1303 4999
rect 2471 4965 2487 4999
rect 1287 4918 2487 4965
rect -2487 71 -1287 118
rect -2487 37 -2471 71
rect -1303 37 -1287 71
rect -2487 21 -1287 37
rect -1229 71 -29 118
rect -1229 37 -1213 71
rect -45 37 -29 71
rect -1229 21 -29 37
rect 29 71 1229 118
rect 29 37 45 71
rect 1213 37 1229 71
rect 29 21 1229 37
rect 1287 71 2487 118
rect 1287 37 1303 71
rect 2471 37 2487 71
rect 1287 21 2487 37
rect -2487 -37 -1287 -21
rect -2487 -71 -2471 -37
rect -1303 -71 -1287 -37
rect -2487 -118 -1287 -71
rect -1229 -37 -29 -21
rect -1229 -71 -1213 -37
rect -45 -71 -29 -37
rect -1229 -118 -29 -71
rect 29 -37 1229 -21
rect 29 -71 45 -37
rect 1213 -71 1229 -37
rect 29 -118 1229 -71
rect 1287 -37 2487 -21
rect 1287 -71 1303 -37
rect 2471 -71 2487 -37
rect 1287 -118 2487 -71
rect -2487 -4965 -1287 -4918
rect -2487 -4999 -2471 -4965
rect -1303 -4999 -1287 -4965
rect -2487 -5015 -1287 -4999
rect -1229 -4965 -29 -4918
rect -1229 -4999 -1213 -4965
rect -45 -4999 -29 -4965
rect -1229 -5015 -29 -4999
rect 29 -4965 1229 -4918
rect 29 -4999 45 -4965
rect 1213 -4999 1229 -4965
rect 29 -5015 1229 -4999
rect 1287 -4965 2487 -4918
rect 1287 -4999 1303 -4965
rect 2471 -4999 2487 -4965
rect 1287 -5015 2487 -4999
rect -2487 -5073 -1287 -5057
rect -2487 -5107 -2471 -5073
rect -1303 -5107 -1287 -5073
rect -2487 -5154 -1287 -5107
rect -1229 -5073 -29 -5057
rect -1229 -5107 -1213 -5073
rect -45 -5107 -29 -5073
rect -1229 -5154 -29 -5107
rect 29 -5073 1229 -5057
rect 29 -5107 45 -5073
rect 1213 -5107 1229 -5073
rect 29 -5154 1229 -5107
rect 1287 -5073 2487 -5057
rect 1287 -5107 1303 -5073
rect 2471 -5107 2487 -5073
rect 1287 -5154 2487 -5107
rect -2487 -10001 -1287 -9954
rect -2487 -10035 -2471 -10001
rect -1303 -10035 -1287 -10001
rect -2487 -10051 -1287 -10035
rect -1229 -10001 -29 -9954
rect -1229 -10035 -1213 -10001
rect -45 -10035 -29 -10001
rect -1229 -10051 -29 -10035
rect 29 -10001 1229 -9954
rect 29 -10035 45 -10001
rect 1213 -10035 1229 -10001
rect 29 -10051 1229 -10035
rect 1287 -10001 2487 -9954
rect 1287 -10035 1303 -10001
rect 2471 -10035 2487 -10001
rect 1287 -10051 2487 -10035
<< polycont >>
rect -2471 10001 -1303 10035
rect -1213 10001 -45 10035
rect 45 10001 1213 10035
rect 1303 10001 2471 10035
rect -2471 5073 -1303 5107
rect -1213 5073 -45 5107
rect 45 5073 1213 5107
rect 1303 5073 2471 5107
rect -2471 4965 -1303 4999
rect -1213 4965 -45 4999
rect 45 4965 1213 4999
rect 1303 4965 2471 4999
rect -2471 37 -1303 71
rect -1213 37 -45 71
rect 45 37 1213 71
rect 1303 37 2471 71
rect -2471 -71 -1303 -37
rect -1213 -71 -45 -37
rect 45 -71 1213 -37
rect 1303 -71 2471 -37
rect -2471 -4999 -1303 -4965
rect -1213 -4999 -45 -4965
rect 45 -4999 1213 -4965
rect 1303 -4999 2471 -4965
rect -2471 -5107 -1303 -5073
rect -1213 -5107 -45 -5073
rect 45 -5107 1213 -5073
rect 1303 -5107 2471 -5073
rect -2471 -10035 -1303 -10001
rect -1213 -10035 -45 -10001
rect 45 -10035 1213 -10001
rect 1303 -10035 2471 -10001
<< locali >>
rect -2667 10139 -2571 10173
rect 2571 10139 2667 10173
rect -2667 10077 -2633 10139
rect 2633 10077 2667 10139
rect -2487 10001 -2471 10035
rect -1303 10001 -1287 10035
rect -1229 10001 -1213 10035
rect -45 10001 -29 10035
rect 29 10001 45 10035
rect 1213 10001 1229 10035
rect 1287 10001 1303 10035
rect 2471 10001 2487 10035
rect -2533 9942 -2499 9958
rect -2533 5150 -2499 5166
rect -1275 9942 -1241 9958
rect -1275 5150 -1241 5166
rect -17 9942 17 9958
rect -17 5150 17 5166
rect 1241 9942 1275 9958
rect 1241 5150 1275 5166
rect 2499 9942 2533 9958
rect 2499 5150 2533 5166
rect -2487 5073 -2471 5107
rect -1303 5073 -1287 5107
rect -1229 5073 -1213 5107
rect -45 5073 -29 5107
rect 29 5073 45 5107
rect 1213 5073 1229 5107
rect 1287 5073 1303 5107
rect 2471 5073 2487 5107
rect -2487 4965 -2471 4999
rect -1303 4965 -1287 4999
rect -1229 4965 -1213 4999
rect -45 4965 -29 4999
rect 29 4965 45 4999
rect 1213 4965 1229 4999
rect 1287 4965 1303 4999
rect 2471 4965 2487 4999
rect -2533 4906 -2499 4922
rect -2533 114 -2499 130
rect -1275 4906 -1241 4922
rect -1275 114 -1241 130
rect -17 4906 17 4922
rect -17 114 17 130
rect 1241 4906 1275 4922
rect 1241 114 1275 130
rect 2499 4906 2533 4922
rect 2499 114 2533 130
rect -2487 37 -2471 71
rect -1303 37 -1287 71
rect -1229 37 -1213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 1213 37 1229 71
rect 1287 37 1303 71
rect 2471 37 2487 71
rect -2487 -71 -2471 -37
rect -1303 -71 -1287 -37
rect -1229 -71 -1213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 1213 -71 1229 -37
rect 1287 -71 1303 -37
rect 2471 -71 2487 -37
rect -2533 -130 -2499 -114
rect -2533 -4922 -2499 -4906
rect -1275 -130 -1241 -114
rect -1275 -4922 -1241 -4906
rect -17 -130 17 -114
rect -17 -4922 17 -4906
rect 1241 -130 1275 -114
rect 1241 -4922 1275 -4906
rect 2499 -130 2533 -114
rect 2499 -4922 2533 -4906
rect -2487 -4999 -2471 -4965
rect -1303 -4999 -1287 -4965
rect -1229 -4999 -1213 -4965
rect -45 -4999 -29 -4965
rect 29 -4999 45 -4965
rect 1213 -4999 1229 -4965
rect 1287 -4999 1303 -4965
rect 2471 -4999 2487 -4965
rect -2487 -5107 -2471 -5073
rect -1303 -5107 -1287 -5073
rect -1229 -5107 -1213 -5073
rect -45 -5107 -29 -5073
rect 29 -5107 45 -5073
rect 1213 -5107 1229 -5073
rect 1287 -5107 1303 -5073
rect 2471 -5107 2487 -5073
rect -2533 -5166 -2499 -5150
rect -2533 -9958 -2499 -9942
rect -1275 -5166 -1241 -5150
rect -1275 -9958 -1241 -9942
rect -17 -5166 17 -5150
rect -17 -9958 17 -9942
rect 1241 -5166 1275 -5150
rect 1241 -9958 1275 -9942
rect 2499 -5166 2533 -5150
rect 2499 -9958 2533 -9942
rect -2487 -10035 -2471 -10001
rect -1303 -10035 -1287 -10001
rect -1229 -10035 -1213 -10001
rect -45 -10035 -29 -10001
rect 29 -10035 45 -10001
rect 1213 -10035 1229 -10001
rect 1287 -10035 1303 -10001
rect 2471 -10035 2487 -10001
rect -2667 -10139 -2633 -10077
rect 2633 -10139 2667 -10077
rect -2667 -10173 -2571 -10139
rect 2571 -10173 2667 -10139
<< viali >>
rect -2471 10001 -1303 10035
rect -1213 10001 -45 10035
rect 45 10001 1213 10035
rect 1303 10001 2471 10035
rect -2533 5166 -2499 9942
rect -1275 5166 -1241 9942
rect -17 5166 17 9942
rect 1241 5166 1275 9942
rect 2499 5166 2533 9942
rect -2471 5073 -1303 5107
rect -1213 5073 -45 5107
rect 45 5073 1213 5107
rect 1303 5073 2471 5107
rect -2471 4965 -1303 4999
rect -1213 4965 -45 4999
rect 45 4965 1213 4999
rect 1303 4965 2471 4999
rect -2533 130 -2499 4906
rect -1275 130 -1241 4906
rect -17 130 17 4906
rect 1241 130 1275 4906
rect 2499 130 2533 4906
rect -2471 37 -1303 71
rect -1213 37 -45 71
rect 45 37 1213 71
rect 1303 37 2471 71
rect -2471 -71 -1303 -37
rect -1213 -71 -45 -37
rect 45 -71 1213 -37
rect 1303 -71 2471 -37
rect -2533 -4906 -2499 -130
rect -1275 -4906 -1241 -130
rect -17 -4906 17 -130
rect 1241 -4906 1275 -130
rect 2499 -4906 2533 -130
rect -2471 -4999 -1303 -4965
rect -1213 -4999 -45 -4965
rect 45 -4999 1213 -4965
rect 1303 -4999 2471 -4965
rect -2471 -5107 -1303 -5073
rect -1213 -5107 -45 -5073
rect 45 -5107 1213 -5073
rect 1303 -5107 2471 -5073
rect -2533 -9942 -2499 -5166
rect -1275 -9942 -1241 -5166
rect -17 -9942 17 -5166
rect 1241 -9942 1275 -5166
rect 2499 -9942 2533 -5166
rect -2471 -10035 -1303 -10001
rect -1213 -10035 -45 -10001
rect 45 -10035 1213 -10001
rect 1303 -10035 2471 -10001
<< metal1 >>
rect -2483 10035 -1291 10041
rect -2483 10001 -2471 10035
rect -1303 10001 -1291 10035
rect -2483 9995 -1291 10001
rect -1225 10035 -33 10041
rect -1225 10001 -1213 10035
rect -45 10001 -33 10035
rect -1225 9995 -33 10001
rect 33 10035 1225 10041
rect 33 10001 45 10035
rect 1213 10001 1225 10035
rect 33 9995 1225 10001
rect 1291 10035 2483 10041
rect 1291 10001 1303 10035
rect 2471 10001 2483 10035
rect 1291 9995 2483 10001
rect -2539 9942 -2493 9954
rect -2539 5166 -2533 9942
rect -2499 5166 -2493 9942
rect -2539 5154 -2493 5166
rect -1281 9942 -1235 9954
rect -1281 5166 -1275 9942
rect -1241 5166 -1235 9942
rect -1281 5154 -1235 5166
rect -23 9942 23 9954
rect -23 5166 -17 9942
rect 17 5166 23 9942
rect -23 5154 23 5166
rect 1235 9942 1281 9954
rect 1235 5166 1241 9942
rect 1275 5166 1281 9942
rect 1235 5154 1281 5166
rect 2493 9942 2539 9954
rect 2493 5166 2499 9942
rect 2533 5166 2539 9942
rect 2493 5154 2539 5166
rect -2483 5107 -1291 5113
rect -2483 5073 -2471 5107
rect -1303 5073 -1291 5107
rect -2483 5067 -1291 5073
rect -1225 5107 -33 5113
rect -1225 5073 -1213 5107
rect -45 5073 -33 5107
rect -1225 5067 -33 5073
rect 33 5107 1225 5113
rect 33 5073 45 5107
rect 1213 5073 1225 5107
rect 33 5067 1225 5073
rect 1291 5107 2483 5113
rect 1291 5073 1303 5107
rect 2471 5073 2483 5107
rect 1291 5067 2483 5073
rect -2483 4999 -1291 5005
rect -2483 4965 -2471 4999
rect -1303 4965 -1291 4999
rect -2483 4959 -1291 4965
rect -1225 4999 -33 5005
rect -1225 4965 -1213 4999
rect -45 4965 -33 4999
rect -1225 4959 -33 4965
rect 33 4999 1225 5005
rect 33 4965 45 4999
rect 1213 4965 1225 4999
rect 33 4959 1225 4965
rect 1291 4999 2483 5005
rect 1291 4965 1303 4999
rect 2471 4965 2483 4999
rect 1291 4959 2483 4965
rect -2539 4906 -2493 4918
rect -2539 130 -2533 4906
rect -2499 130 -2493 4906
rect -2539 118 -2493 130
rect -1281 4906 -1235 4918
rect -1281 130 -1275 4906
rect -1241 130 -1235 4906
rect -1281 118 -1235 130
rect -23 4906 23 4918
rect -23 130 -17 4906
rect 17 130 23 4906
rect -23 118 23 130
rect 1235 4906 1281 4918
rect 1235 130 1241 4906
rect 1275 130 1281 4906
rect 1235 118 1281 130
rect 2493 4906 2539 4918
rect 2493 130 2499 4906
rect 2533 130 2539 4906
rect 2493 118 2539 130
rect -2483 71 -1291 77
rect -2483 37 -2471 71
rect -1303 37 -1291 71
rect -2483 31 -1291 37
rect -1225 71 -33 77
rect -1225 37 -1213 71
rect -45 37 -33 71
rect -1225 31 -33 37
rect 33 71 1225 77
rect 33 37 45 71
rect 1213 37 1225 71
rect 33 31 1225 37
rect 1291 71 2483 77
rect 1291 37 1303 71
rect 2471 37 2483 71
rect 1291 31 2483 37
rect -2483 -37 -1291 -31
rect -2483 -71 -2471 -37
rect -1303 -71 -1291 -37
rect -2483 -77 -1291 -71
rect -1225 -37 -33 -31
rect -1225 -71 -1213 -37
rect -45 -71 -33 -37
rect -1225 -77 -33 -71
rect 33 -37 1225 -31
rect 33 -71 45 -37
rect 1213 -71 1225 -37
rect 33 -77 1225 -71
rect 1291 -37 2483 -31
rect 1291 -71 1303 -37
rect 2471 -71 2483 -37
rect 1291 -77 2483 -71
rect -2539 -130 -2493 -118
rect -2539 -4906 -2533 -130
rect -2499 -4906 -2493 -130
rect -2539 -4918 -2493 -4906
rect -1281 -130 -1235 -118
rect -1281 -4906 -1275 -130
rect -1241 -4906 -1235 -130
rect -1281 -4918 -1235 -4906
rect -23 -130 23 -118
rect -23 -4906 -17 -130
rect 17 -4906 23 -130
rect -23 -4918 23 -4906
rect 1235 -130 1281 -118
rect 1235 -4906 1241 -130
rect 1275 -4906 1281 -130
rect 1235 -4918 1281 -4906
rect 2493 -130 2539 -118
rect 2493 -4906 2499 -130
rect 2533 -4906 2539 -130
rect 2493 -4918 2539 -4906
rect -2483 -4965 -1291 -4959
rect -2483 -4999 -2471 -4965
rect -1303 -4999 -1291 -4965
rect -2483 -5005 -1291 -4999
rect -1225 -4965 -33 -4959
rect -1225 -4999 -1213 -4965
rect -45 -4999 -33 -4965
rect -1225 -5005 -33 -4999
rect 33 -4965 1225 -4959
rect 33 -4999 45 -4965
rect 1213 -4999 1225 -4965
rect 33 -5005 1225 -4999
rect 1291 -4965 2483 -4959
rect 1291 -4999 1303 -4965
rect 2471 -4999 2483 -4965
rect 1291 -5005 2483 -4999
rect -2483 -5073 -1291 -5067
rect -2483 -5107 -2471 -5073
rect -1303 -5107 -1291 -5073
rect -2483 -5113 -1291 -5107
rect -1225 -5073 -33 -5067
rect -1225 -5107 -1213 -5073
rect -45 -5107 -33 -5073
rect -1225 -5113 -33 -5107
rect 33 -5073 1225 -5067
rect 33 -5107 45 -5073
rect 1213 -5107 1225 -5073
rect 33 -5113 1225 -5107
rect 1291 -5073 2483 -5067
rect 1291 -5107 1303 -5073
rect 2471 -5107 2483 -5073
rect 1291 -5113 2483 -5107
rect -2539 -5166 -2493 -5154
rect -2539 -9942 -2533 -5166
rect -2499 -9942 -2493 -5166
rect -2539 -9954 -2493 -9942
rect -1281 -5166 -1235 -5154
rect -1281 -9942 -1275 -5166
rect -1241 -9942 -1235 -5166
rect -1281 -9954 -1235 -9942
rect -23 -5166 23 -5154
rect -23 -9942 -17 -5166
rect 17 -9942 23 -5166
rect -23 -9954 23 -9942
rect 1235 -5166 1281 -5154
rect 1235 -9942 1241 -5166
rect 1275 -9942 1281 -5166
rect 1235 -9954 1281 -9942
rect 2493 -5166 2539 -5154
rect 2493 -9942 2499 -5166
rect 2533 -9942 2539 -5166
rect 2493 -9954 2539 -9942
rect -2483 -10001 -1291 -9995
rect -2483 -10035 -2471 -10001
rect -1303 -10035 -1291 -10001
rect -2483 -10041 -1291 -10035
rect -1225 -10001 -33 -9995
rect -1225 -10035 -1213 -10001
rect -45 -10035 -33 -10001
rect -1225 -10041 -33 -10035
rect 33 -10001 1225 -9995
rect 33 -10035 45 -10001
rect 1213 -10035 1225 -10001
rect 33 -10041 1225 -10035
rect 1291 -10001 2483 -9995
rect 1291 -10035 1303 -10001
rect 2471 -10035 2483 -10001
rect 1291 -10041 2483 -10035
<< properties >>
string FIXED_BBOX -2650 -10156 2650 10156
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 24.0 l 6.0 m 4 nf 4 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
