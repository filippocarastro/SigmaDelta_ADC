magic
tech sky130B
magscale 1 2
timestamp 1667069721
<< nwell >>
rect -858 -20087 858 20087
<< mvpmos >>
rect -600 13390 600 19790
rect -600 6754 600 13154
rect -600 118 600 6518
rect -600 -6518 600 -118
rect -600 -13154 600 -6754
rect -600 -19790 600 -13390
<< mvpdiff >>
rect -658 19778 -600 19790
rect -658 13402 -646 19778
rect -612 13402 -600 19778
rect -658 13390 -600 13402
rect 600 19778 658 19790
rect 600 13402 612 19778
rect 646 13402 658 19778
rect 600 13390 658 13402
rect -658 13142 -600 13154
rect -658 6766 -646 13142
rect -612 6766 -600 13142
rect -658 6754 -600 6766
rect 600 13142 658 13154
rect 600 6766 612 13142
rect 646 6766 658 13142
rect 600 6754 658 6766
rect -658 6506 -600 6518
rect -658 130 -646 6506
rect -612 130 -600 6506
rect -658 118 -600 130
rect 600 6506 658 6518
rect 600 130 612 6506
rect 646 130 658 6506
rect 600 118 658 130
rect -658 -130 -600 -118
rect -658 -6506 -646 -130
rect -612 -6506 -600 -130
rect -658 -6518 -600 -6506
rect 600 -130 658 -118
rect 600 -6506 612 -130
rect 646 -6506 658 -130
rect 600 -6518 658 -6506
rect -658 -6766 -600 -6754
rect -658 -13142 -646 -6766
rect -612 -13142 -600 -6766
rect -658 -13154 -600 -13142
rect 600 -6766 658 -6754
rect 600 -13142 612 -6766
rect 646 -13142 658 -6766
rect 600 -13154 658 -13142
rect -658 -13402 -600 -13390
rect -658 -19778 -646 -13402
rect -612 -19778 -600 -13402
rect -658 -19790 -600 -19778
rect 600 -13402 658 -13390
rect 600 -19778 612 -13402
rect 646 -19778 658 -13402
rect 600 -19790 658 -19778
<< mvpdiffc >>
rect -646 13402 -612 19778
rect 612 13402 646 19778
rect -646 6766 -612 13142
rect 612 6766 646 13142
rect -646 130 -612 6506
rect 612 130 646 6506
rect -646 -6506 -612 -130
rect 612 -6506 646 -130
rect -646 -13142 -612 -6766
rect 612 -13142 646 -6766
rect -646 -19778 -612 -13402
rect 612 -19778 646 -13402
<< mvnsubdiff >>
rect -792 20009 792 20021
rect -792 19975 -684 20009
rect 684 19975 792 20009
rect -792 19963 792 19975
rect -792 19913 -734 19963
rect -792 -19913 -780 19913
rect -746 -19913 -734 19913
rect 734 19913 792 19963
rect -792 -19963 -734 -19913
rect 734 -19913 746 19913
rect 780 -19913 792 19913
rect 734 -19963 792 -19913
rect -792 -19975 792 -19963
rect -792 -20009 -684 -19975
rect 684 -20009 792 -19975
rect -792 -20021 792 -20009
<< mvnsubdiffcont >>
rect -684 19975 684 20009
rect -780 -19913 -746 19913
rect 746 -19913 780 19913
rect -684 -20009 684 -19975
<< poly >>
rect -600 19871 600 19887
rect -600 19837 -584 19871
rect 584 19837 600 19871
rect -600 19790 600 19837
rect -600 13343 600 13390
rect -600 13309 -584 13343
rect 584 13309 600 13343
rect -600 13293 600 13309
rect -600 13235 600 13251
rect -600 13201 -584 13235
rect 584 13201 600 13235
rect -600 13154 600 13201
rect -600 6707 600 6754
rect -600 6673 -584 6707
rect 584 6673 600 6707
rect -600 6657 600 6673
rect -600 6599 600 6615
rect -600 6565 -584 6599
rect 584 6565 600 6599
rect -600 6518 600 6565
rect -600 71 600 118
rect -600 37 -584 71
rect 584 37 600 71
rect -600 21 600 37
rect -600 -37 600 -21
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -600 -118 600 -71
rect -600 -6565 600 -6518
rect -600 -6599 -584 -6565
rect 584 -6599 600 -6565
rect -600 -6615 600 -6599
rect -600 -6673 600 -6657
rect -600 -6707 -584 -6673
rect 584 -6707 600 -6673
rect -600 -6754 600 -6707
rect -600 -13201 600 -13154
rect -600 -13235 -584 -13201
rect 584 -13235 600 -13201
rect -600 -13251 600 -13235
rect -600 -13309 600 -13293
rect -600 -13343 -584 -13309
rect 584 -13343 600 -13309
rect -600 -13390 600 -13343
rect -600 -19837 600 -19790
rect -600 -19871 -584 -19837
rect 584 -19871 600 -19837
rect -600 -19887 600 -19871
<< polycont >>
rect -584 19837 584 19871
rect -584 13309 584 13343
rect -584 13201 584 13235
rect -584 6673 584 6707
rect -584 6565 584 6599
rect -584 37 584 71
rect -584 -71 584 -37
rect -584 -6599 584 -6565
rect -584 -6707 584 -6673
rect -584 -13235 584 -13201
rect -584 -13343 584 -13309
rect -584 -19871 584 -19837
<< locali >>
rect -780 19975 -684 20009
rect 684 19975 780 20009
rect -780 19913 -746 19975
rect 746 19913 780 19975
rect -600 19837 -584 19871
rect 584 19837 600 19871
rect -646 19778 -612 19794
rect -646 13386 -612 13402
rect 612 19778 646 19794
rect 612 13386 646 13402
rect -600 13309 -584 13343
rect 584 13309 600 13343
rect -600 13201 -584 13235
rect 584 13201 600 13235
rect -646 13142 -612 13158
rect -646 6750 -612 6766
rect 612 13142 646 13158
rect 612 6750 646 6766
rect -600 6673 -584 6707
rect 584 6673 600 6707
rect -600 6565 -584 6599
rect 584 6565 600 6599
rect -646 6506 -612 6522
rect -646 114 -612 130
rect 612 6506 646 6522
rect 612 114 646 130
rect -600 37 -584 71
rect 584 37 600 71
rect -600 -71 -584 -37
rect 584 -71 600 -37
rect -646 -130 -612 -114
rect -646 -6522 -612 -6506
rect 612 -130 646 -114
rect 612 -6522 646 -6506
rect -600 -6599 -584 -6565
rect 584 -6599 600 -6565
rect -600 -6707 -584 -6673
rect 584 -6707 600 -6673
rect -646 -6766 -612 -6750
rect -646 -13158 -612 -13142
rect 612 -6766 646 -6750
rect 612 -13158 646 -13142
rect -600 -13235 -584 -13201
rect 584 -13235 600 -13201
rect -600 -13343 -584 -13309
rect 584 -13343 600 -13309
rect -646 -13402 -612 -13386
rect -646 -19794 -612 -19778
rect 612 -13402 646 -13386
rect 612 -19794 646 -19778
rect -600 -19871 -584 -19837
rect 584 -19871 600 -19837
rect -780 -19975 -746 -19913
rect 746 -19975 780 -19913
rect -780 -20009 -684 -19975
rect 684 -20009 780 -19975
<< viali >>
rect -584 19837 584 19871
rect -646 13402 -612 19778
rect 612 13402 646 19778
rect -584 13309 584 13343
rect -584 13201 584 13235
rect -646 6766 -612 13142
rect 612 6766 646 13142
rect -584 6673 584 6707
rect -584 6565 584 6599
rect -646 130 -612 6506
rect 612 130 646 6506
rect -584 37 584 71
rect -584 -71 584 -37
rect -646 -6506 -612 -130
rect 612 -6506 646 -130
rect -584 -6599 584 -6565
rect -584 -6707 584 -6673
rect -646 -13142 -612 -6766
rect 612 -13142 646 -6766
rect -584 -13235 584 -13201
rect -584 -13343 584 -13309
rect -646 -19778 -612 -13402
rect 612 -19778 646 -13402
rect -584 -19871 584 -19837
<< metal1 >>
rect -596 19871 596 19877
rect -596 19837 -584 19871
rect 584 19837 596 19871
rect -596 19831 596 19837
rect -652 19778 -606 19790
rect -652 13402 -646 19778
rect -612 13402 -606 19778
rect -652 13390 -606 13402
rect 606 19778 652 19790
rect 606 13402 612 19778
rect 646 13402 652 19778
rect 606 13390 652 13402
rect -596 13343 596 13349
rect -596 13309 -584 13343
rect 584 13309 596 13343
rect -596 13303 596 13309
rect -596 13235 596 13241
rect -596 13201 -584 13235
rect 584 13201 596 13235
rect -596 13195 596 13201
rect -652 13142 -606 13154
rect -652 6766 -646 13142
rect -612 6766 -606 13142
rect -652 6754 -606 6766
rect 606 13142 652 13154
rect 606 6766 612 13142
rect 646 6766 652 13142
rect 606 6754 652 6766
rect -596 6707 596 6713
rect -596 6673 -584 6707
rect 584 6673 596 6707
rect -596 6667 596 6673
rect -596 6599 596 6605
rect -596 6565 -584 6599
rect 584 6565 596 6599
rect -596 6559 596 6565
rect -652 6506 -606 6518
rect -652 130 -646 6506
rect -612 130 -606 6506
rect -652 118 -606 130
rect 606 6506 652 6518
rect 606 130 612 6506
rect 646 130 652 6506
rect 606 118 652 130
rect -596 71 596 77
rect -596 37 -584 71
rect 584 37 596 71
rect -596 31 596 37
rect -596 -37 596 -31
rect -596 -71 -584 -37
rect 584 -71 596 -37
rect -596 -77 596 -71
rect -652 -130 -606 -118
rect -652 -6506 -646 -130
rect -612 -6506 -606 -130
rect -652 -6518 -606 -6506
rect 606 -130 652 -118
rect 606 -6506 612 -130
rect 646 -6506 652 -130
rect 606 -6518 652 -6506
rect -596 -6565 596 -6559
rect -596 -6599 -584 -6565
rect 584 -6599 596 -6565
rect -596 -6605 596 -6599
rect -596 -6673 596 -6667
rect -596 -6707 -584 -6673
rect 584 -6707 596 -6673
rect -596 -6713 596 -6707
rect -652 -6766 -606 -6754
rect -652 -13142 -646 -6766
rect -612 -13142 -606 -6766
rect -652 -13154 -606 -13142
rect 606 -6766 652 -6754
rect 606 -13142 612 -6766
rect 646 -13142 652 -6766
rect 606 -13154 652 -13142
rect -596 -13201 596 -13195
rect -596 -13235 -584 -13201
rect 584 -13235 596 -13201
rect -596 -13241 596 -13235
rect -596 -13309 596 -13303
rect -596 -13343 -584 -13309
rect 584 -13343 596 -13309
rect -596 -13349 596 -13343
rect -652 -13402 -606 -13390
rect -652 -19778 -646 -13402
rect -612 -19778 -606 -13402
rect -652 -19790 -606 -19778
rect 606 -13402 652 -13390
rect 606 -19778 612 -13402
rect 646 -19778 652 -13402
rect 606 -19790 652 -19778
rect -596 -19837 596 -19831
rect -596 -19871 -584 -19837
rect 584 -19871 596 -19837
rect -596 -19877 596 -19871
<< properties >>
string FIXED_BBOX -763 -19992 763 19992
string gencell sky130_fd_pr__pfet_g5v0d10v5
string library sky130
string parameters w 32.0 l 6.0 m 6 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.50 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
