VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OpAmp
  CLASS BLOCK ;
  FOREIGN OpAmp ;
  ORIGIN -58.760 -69.940 ;
  SIZE 168.280 BY 113.250 ;
  PIN Vinn
    PORT
      LAYER met1 ;
        RECT 133.020 140.460 140.020 142.490 ;
    END
  END Vinn
  PIN Vinp
    PORT
      LAYER met1 ;
        RECT 218.950 140.950 227.040 143.010 ;
    END
  END Vinp
  PIN GND
    PORT
      LAYER met1 ;
        RECT 58.760 69.940 226.110 80.070 ;
    END
  END GND
  PIN VDD
    PORT
      LAYER met1 ;
        RECT 59.940 175.510 210.020 183.190 ;
    END
  END VDD
  PIN Ibias
    PORT
      LAYER met1 ;
        RECT 74.175 147.495 226.645 149.005 ;
    END
  END Ibias
  PIN Vout
    PORT
      LAYER met1 ;
        RECT 69.240 140.140 70.240 141.140 ;
    END
  END Vout
  OBS
      LAYER li1 ;
        RECT 69.530 79.490 220.560 176.400 ;
      LAYER met1 ;
        RECT 58.760 175.230 59.660 183.190 ;
        RECT 210.300 175.230 226.880 183.190 ;
        RECT 58.760 149.285 226.880 175.230 ;
        RECT 58.760 147.215 73.895 149.285 ;
        RECT 58.760 143.290 226.880 147.215 ;
        RECT 58.760 142.770 218.670 143.290 ;
        RECT 58.760 141.420 132.740 142.770 ;
        RECT 58.760 139.860 68.960 141.420 ;
        RECT 70.520 140.180 132.740 141.420 ;
        RECT 140.300 140.670 218.670 142.770 ;
        RECT 140.300 140.180 226.880 140.670 ;
        RECT 70.520 139.860 226.880 140.180 ;
        RECT 58.760 80.350 226.880 139.860 ;
        RECT 58.760 80.070 219.150 80.180 ;
        RECT 226.390 80.070 226.880 80.350 ;
      LAYER met2 ;
        RECT 67.800 81.990 226.850 174.970 ;
      LAYER met3 ;
        RECT 104.700 86.500 136.195 121.495 ;
      LAYER met4 ;
        RECT 105.395 86.560 136.175 117.440 ;
  END
END OpAmp
END LIBRARY

